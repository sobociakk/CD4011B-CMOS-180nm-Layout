magic
tech scmos
timestamp 1769391498
<< metal1 >>
rect 6846 3052 7546 3239
rect 6846 2837 7614 3052
rect 6846 2639 7546 2837
<< metal2 >>
rect 6512 4411 6520 4414
rect 6846 2639 7546 3239
rect 9186 1667 9189 1675
<< metal3 >>
rect 6846 2639 7546 3239
<< metal4 >>
rect 6846 2639 7546 3239
<< m6contact >>
rect 6846 2639 7546 3239
<< glass >>
rect 6876 2669 7516 3209
<< end >>
