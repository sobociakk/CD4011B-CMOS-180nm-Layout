magic
tech scmos
timestamp 1769746565
<< nwell >>
rect -5104 226 -4856 323
rect -5208 130 -4856 226
rect -5286 94 -4856 130
rect -5269 86 -4856 94
rect -5269 74 -5202 86
rect -4874 81 -4856 86
<< ntransistor >>
rect -5258 63 -5256 66
rect -5239 63 -5237 66
rect -5215 63 -5213 66
rect -5185 49 -5183 52
rect -5254 34 -5252 37
rect -5237 34 -5235 37
rect -5160 26 -5158 53
rect -5136 26 -5134 53
rect -5128 26 -5126 53
rect -5120 26 -5118 53
rect -5112 26 -5110 53
rect -5104 26 -5102 53
rect -5096 26 -5094 53
rect -5088 26 -5086 53
rect -5080 26 -5078 53
rect -5072 26 -5070 53
rect -5049 -47 -5047 53
rect -5041 -47 -5039 53
rect -5033 -47 -5031 53
rect -5025 -47 -5023 53
rect -5017 -47 -5015 53
rect -5009 -47 -5007 53
rect -5001 -47 -4999 53
rect -4993 -47 -4991 53
rect -4985 -47 -4983 53
rect -4977 -47 -4975 53
rect -4969 -47 -4967 53
rect -4961 -47 -4959 53
rect -4953 -47 -4951 53
rect -4945 -47 -4943 53
rect -4937 -47 -4935 53
rect -4929 -47 -4927 53
rect -4921 -47 -4919 53
rect -4913 -47 -4911 53
rect -4905 -47 -4903 53
rect -4897 -47 -4895 53
rect -4889 -47 -4887 53
rect -4881 -47 -4879 53
<< ptransistor >>
rect -5258 101 -5256 107
rect -5250 101 -5248 107
rect -5185 92 -5183 98
rect -5160 92 -5158 146
rect -5136 92 -5134 146
rect -5128 92 -5126 146
rect -5120 92 -5118 146
rect -5112 92 -5110 146
rect -5104 92 -5102 146
rect -5096 92 -5094 146
rect -5088 92 -5086 146
rect -5080 92 -5078 146
rect -5072 92 -5070 146
rect -5049 92 -5047 292
rect -5041 92 -5039 292
rect -5033 92 -5031 292
rect -5025 92 -5023 292
rect -5017 92 -5015 292
rect -5009 92 -5007 292
rect -5001 92 -4999 292
rect -4993 92 -4991 292
rect -4985 92 -4983 292
rect -4977 92 -4975 292
rect -4969 92 -4967 292
rect -4961 92 -4959 292
rect -4953 92 -4951 292
rect -4945 92 -4943 292
rect -4937 92 -4935 292
rect -4929 92 -4927 292
rect -4921 92 -4919 292
rect -4913 92 -4911 292
rect -4905 92 -4903 292
rect -4897 92 -4895 292
rect -4889 92 -4887 292
rect -4881 92 -4879 292
rect -5258 80 -5256 86
rect -5239 80 -5237 86
rect -5215 80 -5213 86
<< ndiffusion >>
rect -5259 63 -5258 66
rect -5256 63 -5255 66
rect -5240 63 -5239 66
rect -5237 63 -5236 66
rect -5216 63 -5215 66
rect -5213 63 -5212 66
rect -5186 49 -5185 52
rect -5183 49 -5182 52
rect -5259 34 -5254 37
rect -5252 34 -5247 37
rect -5243 34 -5237 37
rect -5235 34 -5226 37
rect -5161 26 -5160 53
rect -5158 26 -5157 53
rect -5137 26 -5136 53
rect -5134 26 -5133 53
rect -5129 26 -5128 53
rect -5126 26 -5125 53
rect -5121 26 -5120 53
rect -5118 26 -5117 53
rect -5113 26 -5112 53
rect -5110 26 -5109 53
rect -5105 26 -5104 53
rect -5102 26 -5101 53
rect -5097 26 -5096 53
rect -5094 26 -5093 53
rect -5089 26 -5088 53
rect -5086 26 -5085 53
rect -5081 26 -5080 53
rect -5078 26 -5077 53
rect -5073 26 -5072 53
rect -5070 26 -5069 53
rect -5050 -47 -5049 53
rect -5047 -47 -5046 53
rect -5042 -47 -5041 53
rect -5039 -47 -5038 53
rect -5034 -47 -5033 53
rect -5031 -47 -5030 53
rect -5026 -47 -5025 53
rect -5023 -47 -5022 53
rect -5018 -47 -5017 53
rect -5015 -47 -5014 53
rect -5010 -47 -5009 53
rect -5007 -47 -5006 53
rect -5002 -47 -5001 53
rect -4999 -47 -4998 53
rect -4994 -47 -4993 53
rect -4991 -47 -4990 53
rect -4986 -47 -4985 53
rect -4983 -47 -4982 53
rect -4978 -47 -4977 53
rect -4975 -47 -4974 53
rect -4970 -47 -4969 53
rect -4967 -47 -4966 53
rect -4962 -47 -4961 53
rect -4959 -47 -4958 53
rect -4954 -47 -4953 53
rect -4951 -47 -4950 53
rect -4946 -47 -4945 53
rect -4943 -47 -4942 53
rect -4938 -47 -4937 53
rect -4935 -47 -4934 53
rect -4930 -47 -4929 53
rect -4927 -47 -4926 53
rect -4922 -47 -4921 53
rect -4919 -47 -4918 53
rect -4914 -47 -4913 53
rect -4911 -47 -4910 53
rect -4906 -47 -4905 53
rect -4903 -47 -4902 53
rect -4898 -47 -4897 53
rect -4895 -47 -4894 53
rect -4890 -47 -4889 53
rect -4887 -47 -4886 53
rect -4882 -47 -4881 53
rect -4879 -47 -4878 53
<< pdiffusion >>
rect -5259 101 -5258 107
rect -5256 101 -5255 107
rect -5251 101 -5250 107
rect -5248 101 -5247 107
rect -5186 92 -5185 98
rect -5183 92 -5182 98
rect -5161 92 -5160 146
rect -5158 92 -5157 146
rect -5137 92 -5136 146
rect -5134 92 -5133 146
rect -5129 92 -5128 146
rect -5126 92 -5125 146
rect -5121 92 -5120 146
rect -5118 92 -5117 146
rect -5113 92 -5112 146
rect -5110 92 -5109 146
rect -5105 92 -5104 146
rect -5102 92 -5101 146
rect -5097 92 -5096 146
rect -5094 92 -5093 146
rect -5089 92 -5088 146
rect -5086 92 -5085 146
rect -5081 92 -5080 146
rect -5078 92 -5077 146
rect -5073 92 -5072 146
rect -5070 92 -5069 146
rect -5050 92 -5049 292
rect -5047 92 -5046 292
rect -5042 92 -5041 292
rect -5039 92 -5038 292
rect -5034 92 -5033 292
rect -5031 92 -5030 292
rect -5026 92 -5025 292
rect -5023 92 -5022 292
rect -5018 92 -5017 292
rect -5015 92 -5014 292
rect -5010 92 -5009 292
rect -5007 92 -5006 292
rect -5002 92 -5001 292
rect -4999 92 -4998 292
rect -4994 92 -4993 292
rect -4991 92 -4990 292
rect -4986 92 -4985 292
rect -4983 92 -4982 292
rect -4978 92 -4977 292
rect -4975 92 -4974 292
rect -4970 92 -4969 292
rect -4967 92 -4966 292
rect -4962 92 -4961 292
rect -4959 92 -4958 292
rect -4954 92 -4953 292
rect -4951 92 -4950 292
rect -4946 92 -4945 292
rect -4943 92 -4942 292
rect -4938 92 -4937 292
rect -4935 92 -4934 292
rect -4930 92 -4929 292
rect -4927 92 -4926 292
rect -4922 92 -4921 292
rect -4919 92 -4918 292
rect -4914 92 -4913 292
rect -4911 92 -4910 292
rect -4906 92 -4905 292
rect -4903 92 -4902 292
rect -4898 92 -4897 292
rect -4895 92 -4894 292
rect -4890 92 -4889 292
rect -4887 92 -4886 292
rect -4882 92 -4881 292
rect -4879 92 -4878 292
rect -5259 80 -5258 86
rect -5256 80 -5255 86
rect -5240 80 -5239 86
rect -5237 80 -5236 86
rect -5216 80 -5215 86
rect -5213 80 -5212 86
<< ndcontact >>
rect -5263 63 -5259 67
rect -5255 63 -5251 67
rect -5244 63 -5240 67
rect -5236 63 -5232 67
rect -5220 63 -5216 67
rect -5212 63 -5208 67
rect -5190 49 -5186 53
rect -5182 49 -5178 53
rect -5263 33 -5259 37
rect -5247 33 -5243 37
rect -5226 33 -5222 37
rect -5165 26 -5161 53
rect -5157 26 -5153 53
rect -5141 26 -5137 53
rect -5133 26 -5129 53
rect -5125 26 -5121 53
rect -5117 26 -5113 53
rect -5109 26 -5105 53
rect -5101 26 -5097 53
rect -5093 26 -5089 53
rect -5085 26 -5081 53
rect -5077 26 -5073 53
rect -5069 26 -5065 53
rect -5054 -47 -5050 53
rect -5046 -47 -5042 53
rect -5038 -47 -5034 53
rect -5030 -47 -5026 53
rect -5022 -47 -5018 53
rect -5014 -47 -5010 53
rect -5006 -47 -5002 53
rect -4998 -47 -4994 53
rect -4990 -47 -4986 53
rect -4982 -47 -4978 53
rect -4974 -47 -4970 53
rect -4966 -47 -4962 53
rect -4958 -47 -4954 53
rect -4950 -47 -4946 53
rect -4942 -47 -4938 53
rect -4934 -47 -4930 53
rect -4926 -47 -4922 53
rect -4918 -47 -4914 53
rect -4910 -47 -4906 53
rect -4902 -47 -4898 53
rect -4894 -47 -4890 53
rect -4886 -47 -4882 53
rect -4878 -47 -4874 53
<< pdcontact >>
rect -5263 101 -5259 107
rect -5255 101 -5251 107
rect -5247 101 -5243 107
rect -5190 92 -5186 98
rect -5182 92 -5178 98
rect -5165 92 -5161 146
rect -5157 92 -5153 146
rect -5141 92 -5137 146
rect -5133 92 -5129 146
rect -5125 92 -5121 146
rect -5117 92 -5113 146
rect -5109 92 -5105 146
rect -5101 92 -5097 146
rect -5093 92 -5089 146
rect -5085 92 -5081 146
rect -5077 92 -5073 146
rect -5069 92 -5065 146
rect -5054 92 -5050 292
rect -5046 92 -5042 292
rect -5038 92 -5034 292
rect -5030 92 -5026 292
rect -5022 92 -5018 292
rect -5014 92 -5010 292
rect -5006 92 -5002 292
rect -4998 92 -4994 292
rect -4990 92 -4986 292
rect -4982 92 -4978 292
rect -4974 92 -4970 292
rect -4966 92 -4962 292
rect -4958 92 -4954 292
rect -4950 92 -4946 292
rect -4942 92 -4938 292
rect -4934 92 -4930 292
rect -4926 92 -4922 292
rect -4918 92 -4914 292
rect -4910 92 -4906 292
rect -4902 92 -4898 292
rect -4894 92 -4890 292
rect -4886 92 -4882 292
rect -4878 92 -4874 292
rect -5263 80 -5259 86
rect -5255 80 -5251 86
rect -5244 80 -5240 86
rect -5236 80 -5232 86
rect -5220 80 -5216 86
rect -5212 80 -5208 86
<< psubstratepdiff >>
rect -5116 332 -4845 334
rect -5116 328 -5105 332
rect -5101 328 -5099 332
rect -5095 328 -5093 332
rect -5089 328 -5087 332
rect -5083 328 -5081 332
rect -5077 328 -5073 332
rect -5069 328 -5067 332
rect -5063 328 -5061 332
rect -5057 328 -5055 332
rect -5051 328 -5049 332
rect -5045 328 -5043 332
rect -5039 328 -5037 332
rect -5033 328 -5031 332
rect -5027 328 -5025 332
rect -5021 328 -5019 332
rect -5015 328 -5013 332
rect -5009 328 -5007 332
rect -5003 328 -4999 332
rect -4995 328 -4993 332
rect -4989 328 -4987 332
rect -4983 328 -4981 332
rect -4977 328 -4975 332
rect -4971 328 -4969 332
rect -4965 328 -4963 332
rect -4959 328 -4957 332
rect -4953 328 -4951 332
rect -4947 328 -4945 332
rect -4941 328 -4939 332
rect -4935 328 -4933 332
rect -4929 328 -4925 332
rect -4921 328 -4919 332
rect -4915 328 -4913 332
rect -4909 328 -4907 332
rect -4903 328 -4901 332
rect -4897 328 -4895 332
rect -4891 328 -4889 332
rect -4885 328 -4883 332
rect -4879 328 -4877 332
rect -4873 328 -4871 332
rect -4867 328 -4865 332
rect -4861 328 -4859 332
rect -4855 328 -4845 332
rect -5116 327 -4845 328
rect -5116 323 -5114 327
rect -5110 326 -4845 327
rect -5110 323 -5108 326
rect -5116 320 -5108 323
rect -4853 322 -4851 326
rect -4847 322 -4845 326
rect -4853 321 -4845 322
rect -5116 316 -5114 320
rect -5110 316 -5108 320
rect -5116 312 -5108 316
rect -5116 308 -5114 312
rect -5110 308 -5108 312
rect -5116 305 -5108 308
rect -5116 301 -5114 305
rect -5110 301 -5108 305
rect -5116 299 -5108 301
rect -5116 295 -5114 299
rect -5110 295 -5108 299
rect -5116 292 -5108 295
rect -5116 288 -5114 292
rect -5110 288 -5108 292
rect -5116 287 -5108 288
rect -5116 283 -5114 287
rect -5110 283 -5108 287
rect -5116 282 -5108 283
rect -5116 278 -5114 282
rect -5110 278 -5108 282
rect -5116 277 -5108 278
rect -5116 273 -5114 277
rect -5110 273 -5108 277
rect -5116 271 -5108 273
rect -5116 267 -5114 271
rect -5110 267 -5108 271
rect -5116 265 -5108 267
rect -5116 261 -5114 265
rect -5110 261 -5108 265
rect -5116 260 -5108 261
rect -5116 256 -5114 260
rect -5110 256 -5108 260
rect -5116 254 -5108 256
rect -5116 250 -5114 254
rect -5110 250 -5108 254
rect -5116 248 -5108 250
rect -5116 244 -5114 248
rect -5110 244 -5108 248
rect -5116 243 -5108 244
rect -5116 239 -5114 243
rect -5110 239 -5108 243
rect -5219 237 -5108 239
rect -5219 233 -5211 237
rect -5207 233 -5205 237
rect -5201 233 -5199 237
rect -5195 233 -5194 237
rect -5190 233 -5139 237
rect -5135 233 -5134 237
rect -5130 233 -5129 237
rect -5125 233 -5122 237
rect -5118 233 -5108 237
rect -5219 231 -5108 233
rect -5219 230 -5211 231
rect -5219 226 -5217 230
rect -5213 226 -5211 230
rect -5219 223 -5211 226
rect -5219 219 -5217 223
rect -5213 219 -5211 223
rect -5219 218 -5211 219
rect -5219 214 -5217 218
rect -5213 214 -5211 218
rect -5219 210 -5211 214
rect -5219 206 -5217 210
rect -5213 206 -5211 210
rect -5219 205 -5211 206
rect -5219 201 -5217 205
rect -5213 201 -5211 205
rect -5219 200 -5211 201
rect -5219 196 -5217 200
rect -5213 196 -5211 200
rect -5219 192 -5211 196
rect -5219 188 -5217 192
rect -5213 188 -5211 192
rect -5219 184 -5211 188
rect -5219 180 -5217 184
rect -5213 180 -5211 184
rect -5219 177 -5211 180
rect -5219 173 -5217 177
rect -5213 173 -5211 177
rect -5219 171 -5211 173
rect -5219 167 -5217 171
rect -5213 167 -5211 171
rect -5219 166 -5211 167
rect -5219 162 -5217 166
rect -5213 162 -5211 166
rect -5219 158 -5211 162
rect -5219 154 -5217 158
rect -5213 154 -5211 158
rect -5219 153 -5211 154
rect -5219 149 -5217 153
rect -5213 149 -5211 153
rect -5219 145 -5211 149
rect -5219 142 -5217 145
rect -5297 141 -5217 142
rect -5213 141 -5211 145
rect -5297 140 -5211 141
rect -5297 136 -5289 140
rect -5285 136 -5283 140
rect -5279 136 -5276 140
rect -5272 136 -5269 140
rect -5265 136 -5262 140
rect -5258 136 -5255 140
rect -5251 136 -5250 140
rect -5246 136 -5245 140
rect -5241 136 -5239 140
rect -5235 136 -5233 140
rect -5229 136 -5227 140
rect -5223 136 -5222 140
rect -5218 136 -5211 140
rect -5297 134 -5211 136
rect -5297 132 -5289 134
rect -5297 128 -5295 132
rect -5291 128 -5289 132
rect -5297 124 -5289 128
rect -5297 120 -5295 124
rect -5291 120 -5289 124
rect -5297 116 -5289 120
rect -5297 112 -5295 116
rect -5291 112 -5289 116
rect -5297 109 -5289 112
rect -5297 105 -5295 109
rect -5291 105 -5289 109
rect -5297 104 -5289 105
rect -5297 100 -5295 104
rect -5291 100 -5289 104
rect -5297 99 -5289 100
rect -5297 95 -5295 99
rect -5291 95 -5289 99
rect -5297 93 -5289 95
rect -5297 89 -5295 93
rect -5291 89 -5289 93
rect -5297 86 -5289 89
rect -5297 82 -5295 86
rect -5291 82 -5289 86
rect -5297 50 -5289 82
rect -4853 317 -4851 321
rect -4847 317 -4845 321
rect -4853 315 -4845 317
rect -4853 311 -4851 315
rect -4847 311 -4845 315
rect -4853 309 -4845 311
rect -4853 305 -4851 309
rect -4847 305 -4845 309
rect -4853 303 -4845 305
rect -4853 299 -4851 303
rect -4847 299 -4845 303
rect -4853 297 -4845 299
rect -4853 293 -4851 297
rect -4847 293 -4845 297
rect -4853 291 -4845 293
rect -4853 287 -4851 291
rect -4847 287 -4845 291
rect -4853 285 -4845 287
rect -4853 281 -4851 285
rect -4847 281 -4845 285
rect -4853 279 -4845 281
rect -4853 275 -4851 279
rect -4847 275 -4845 279
rect -4853 273 -4845 275
rect -4853 269 -4851 273
rect -4847 269 -4845 273
rect -4853 267 -4845 269
rect -4853 263 -4851 267
rect -4847 263 -4845 267
rect -4853 261 -4845 263
rect -4853 257 -4851 261
rect -4847 257 -4845 261
rect -4853 255 -4845 257
rect -4853 251 -4851 255
rect -4847 251 -4845 255
rect -4853 247 -4845 251
rect -4853 243 -4851 247
rect -4847 243 -4845 247
rect -4853 241 -4845 243
rect -4853 237 -4851 241
rect -4847 237 -4845 241
rect -4853 235 -4845 237
rect -4853 231 -4851 235
rect -4847 231 -4845 235
rect -4853 229 -4845 231
rect -4853 225 -4851 229
rect -4847 225 -4845 229
rect -4853 223 -4845 225
rect -4853 219 -4851 223
rect -4847 219 -4845 223
rect -4853 217 -4845 219
rect -4853 213 -4851 217
rect -4847 213 -4845 217
rect -4853 211 -4845 213
rect -4853 207 -4851 211
rect -4847 207 -4845 211
rect -4853 205 -4845 207
rect -4853 201 -4851 205
rect -4847 201 -4845 205
rect -4853 199 -4845 201
rect -4853 195 -4851 199
rect -4847 195 -4845 199
rect -4853 193 -4845 195
rect -4853 189 -4851 193
rect -4847 189 -4845 193
rect -4853 187 -4845 189
rect -4853 183 -4851 187
rect -4847 183 -4845 187
rect -4853 181 -4845 183
rect -4853 177 -4851 181
rect -4847 177 -4845 181
rect -4853 173 -4845 177
rect -4853 169 -4851 173
rect -4847 169 -4845 173
rect -4853 167 -4845 169
rect -4853 163 -4851 167
rect -4847 163 -4845 167
rect -4853 161 -4845 163
rect -4853 157 -4851 161
rect -4847 157 -4845 161
rect -4853 155 -4845 157
rect -4853 151 -4851 155
rect -4847 151 -4845 155
rect -4853 149 -4845 151
rect -4853 145 -4851 149
rect -4847 145 -4845 149
rect -4853 143 -4845 145
rect -4853 139 -4851 143
rect -4847 139 -4845 143
rect -4853 137 -4845 139
rect -4853 133 -4851 137
rect -4847 133 -4845 137
rect -4853 131 -4845 133
rect -4853 127 -4851 131
rect -4847 127 -4845 131
rect -4853 125 -4845 127
rect -4853 121 -4851 125
rect -4847 121 -4845 125
rect -4853 119 -4845 121
rect -4853 115 -4851 119
rect -4847 115 -4845 119
rect -4853 113 -4845 115
rect -4853 109 -4851 113
rect -4847 109 -4845 113
rect -4853 107 -4845 109
rect -4853 103 -4851 107
rect -4847 103 -4845 107
rect -4853 99 -4845 103
rect -4853 95 -4851 99
rect -4847 95 -4845 99
rect -4853 93 -4845 95
rect -4853 89 -4851 93
rect -4847 89 -4845 93
rect -4853 87 -4845 89
rect -5297 46 -5295 50
rect -5291 46 -5289 50
rect -5297 45 -5289 46
rect -5297 41 -5295 45
rect -5291 41 -5289 45
rect -5297 37 -5289 41
rect -4853 83 -4851 87
rect -4847 83 -4845 87
rect -4853 63 -4845 83
rect -4853 59 -4851 63
rect -4847 59 -4845 63
rect -4853 57 -4845 59
rect -4853 53 -4851 57
rect -4847 53 -4845 57
rect -5297 33 -5295 37
rect -5291 33 -5289 37
rect -5297 29 -5289 33
rect -5297 25 -5295 29
rect -5291 25 -5289 29
rect -5297 21 -5289 25
rect -5297 17 -5295 21
rect -5291 17 -5289 21
rect -5297 16 -5289 17
rect -5297 14 -5063 16
rect -5297 10 -5288 14
rect -5284 10 -5281 14
rect -5277 10 -5275 14
rect -5271 10 -5205 14
rect -5201 10 -5197 14
rect -5193 10 -5189 14
rect -5185 10 -5181 14
rect -5177 10 -5173 14
rect -5169 10 -5167 14
rect -5163 10 -5157 14
rect -5153 10 -5149 14
rect -5145 10 -5141 14
rect -5137 10 -5133 14
rect -5129 10 -5124 14
rect -5120 10 -5117 14
rect -5113 10 -5111 14
rect -5107 10 -5106 14
rect -5102 10 -5101 14
rect -5097 10 -5096 14
rect -5092 10 -5091 14
rect -5087 10 -5086 14
rect -5082 10 -5078 14
rect -5074 10 -5063 14
rect -5297 9 -5063 10
rect -5297 8 -5069 9
rect -5071 5 -5069 8
rect -5065 5 -5063 9
rect -5071 2 -5063 5
rect -5071 -2 -5069 2
rect -5065 -2 -5063 2
rect -5071 -4 -5063 -2
rect -5071 -8 -5069 -4
rect -5065 -8 -5063 -4
rect -5071 -9 -5063 -8
rect -5071 -13 -5069 -9
rect -5065 -13 -5063 -9
rect -5071 -16 -5063 -13
rect -5071 -20 -5069 -16
rect -5065 -20 -5063 -16
rect -5071 -24 -5063 -20
rect -5071 -28 -5069 -24
rect -5065 -28 -5063 -24
rect -5071 -31 -5063 -28
rect -5071 -35 -5069 -31
rect -5065 -35 -5063 -31
rect -5071 -37 -5063 -35
rect -5071 -41 -5069 -37
rect -5065 -41 -5063 -37
rect -5071 -44 -5063 -41
rect -5071 -48 -5069 -44
rect -5065 -48 -5063 -44
rect -4853 51 -4845 53
rect -4853 47 -4851 51
rect -4847 47 -4845 51
rect -4853 45 -4845 47
rect -4853 41 -4851 45
rect -4847 41 -4845 45
rect -4853 39 -4845 41
rect -4853 35 -4851 39
rect -4847 35 -4845 39
rect -4853 33 -4845 35
rect -4853 29 -4851 33
rect -4847 29 -4845 33
rect -4853 25 -4845 29
rect -4853 21 -4851 25
rect -4847 21 -4845 25
rect -4853 19 -4845 21
rect -4853 15 -4851 19
rect -4847 15 -4845 19
rect -4853 13 -4845 15
rect -4853 9 -4851 13
rect -4847 9 -4845 13
rect -4853 7 -4845 9
rect -4853 3 -4851 7
rect -4847 3 -4845 7
rect -4853 1 -4845 3
rect -4853 -3 -4851 1
rect -4847 -3 -4845 1
rect -4853 -5 -4845 -3
rect -4853 -9 -4851 -5
rect -4847 -9 -4845 -5
rect -4853 -11 -4845 -9
rect -4853 -15 -4851 -11
rect -4847 -15 -4845 -11
rect -4853 -17 -4845 -15
rect -4853 -21 -4851 -17
rect -4847 -21 -4845 -17
rect -4853 -23 -4845 -21
rect -4853 -27 -4851 -23
rect -4847 -27 -4845 -23
rect -4853 -29 -4845 -27
rect -4853 -33 -4851 -29
rect -4847 -33 -4845 -29
rect -4853 -35 -4845 -33
rect -4853 -39 -4851 -35
rect -4847 -39 -4845 -35
rect -4853 -41 -4845 -39
rect -4853 -45 -4851 -41
rect -4847 -45 -4845 -41
rect -4853 -46 -4845 -45
rect -5071 -51 -5063 -48
rect -4853 -50 -4851 -46
rect -4847 -50 -4845 -46
rect -5071 -55 -5069 -51
rect -5065 -55 -5063 -51
rect -5071 -56 -5063 -55
rect -4853 -52 -4845 -50
rect -4853 -56 -4851 -52
rect -4847 -56 -4845 -52
rect -5071 -58 -4845 -56
rect -5071 -62 -5062 -58
rect -5058 -62 -5056 -58
rect -5052 -62 -5050 -58
rect -5046 -62 -5044 -58
rect -5040 -62 -5038 -58
rect -5034 -62 -5032 -58
rect -5028 -62 -5026 -58
rect -5022 -62 -5020 -58
rect -5016 -62 -5014 -58
rect -5010 -62 -5006 -58
rect -5002 -62 -5000 -58
rect -4996 -62 -4994 -58
rect -4990 -62 -4988 -58
rect -4984 -62 -4982 -58
rect -4978 -62 -4976 -58
rect -4972 -62 -4970 -58
rect -4966 -62 -4964 -58
rect -4960 -62 -4958 -58
rect -4954 -62 -4952 -58
rect -4948 -62 -4946 -58
rect -4942 -62 -4940 -58
rect -4936 -62 -4932 -58
rect -4928 -62 -4926 -58
rect -4922 -62 -4920 -58
rect -4916 -62 -4914 -58
rect -4910 -62 -4908 -58
rect -4904 -62 -4902 -58
rect -4898 -62 -4896 -58
rect -4892 -62 -4890 -58
rect -4886 -62 -4884 -58
rect -4880 -62 -4878 -58
rect -4874 -62 -4872 -58
rect -4868 -62 -4866 -58
rect -4862 -62 -4861 -58
rect -4857 -62 -4856 -58
rect -4852 -62 -4845 -58
rect -5071 -64 -4845 -62
<< nsubstratendiff >>
rect -5097 318 -4860 320
rect -5097 314 -5088 318
rect -5084 314 -5083 318
rect -5079 314 -5078 318
rect -5074 314 -5072 318
rect -5068 314 -5066 318
rect -5062 314 -5058 318
rect -5054 314 -5052 318
rect -5048 314 -5046 318
rect -5042 314 -5040 318
rect -5036 314 -5034 318
rect -5030 314 -5028 318
rect -5024 314 -5022 318
rect -5018 314 -5016 318
rect -5012 314 -5010 318
rect -5006 314 -5004 318
rect -5000 314 -4998 318
rect -4994 314 -4992 318
rect -4988 314 -4986 318
rect -4982 314 -4980 318
rect -4976 314 -4974 318
rect -4970 314 -4968 318
rect -4964 314 -4962 318
rect -4958 314 -4956 318
rect -4952 314 -4950 318
rect -4946 314 -4944 318
rect -4940 314 -4938 318
rect -4934 314 -4932 318
rect -4928 314 -4926 318
rect -4922 314 -4920 318
rect -4916 314 -4914 318
rect -4910 314 -4908 318
rect -4904 314 -4902 318
rect -4898 314 -4896 318
rect -4892 314 -4890 318
rect -4886 314 -4884 318
rect -4880 314 -4878 318
rect -4874 314 -4872 318
rect -4868 314 -4860 318
rect -5097 313 -4866 314
rect -5097 309 -5095 313
rect -5091 312 -4866 313
rect -5091 309 -5089 312
rect -5097 307 -5089 309
rect -5097 303 -5095 307
rect -5091 303 -5089 307
rect -5097 301 -5089 303
rect -5097 297 -5095 301
rect -5091 297 -5089 301
rect -5097 295 -5089 297
rect -4868 310 -4866 312
rect -4862 310 -4860 314
rect -4868 308 -4860 310
rect -4868 304 -4866 308
rect -4862 304 -4860 308
rect -4868 302 -4860 304
rect -4868 298 -4866 302
rect -4862 298 -4860 302
rect -4868 296 -4860 298
rect -5097 291 -5095 295
rect -5091 291 -5089 295
rect -4868 292 -4866 296
rect -4862 292 -4860 296
rect -5097 289 -5089 291
rect -5097 285 -5095 289
rect -5091 285 -5089 289
rect -5097 281 -5089 285
rect -5097 277 -5095 281
rect -5091 277 -5089 281
rect -5097 275 -5089 277
rect -5097 271 -5095 275
rect -5091 271 -5089 275
rect -5097 267 -5089 271
rect -5097 263 -5095 267
rect -5091 263 -5089 267
rect -5097 259 -5089 263
rect -5097 255 -5095 259
rect -5091 255 -5089 259
rect -5097 253 -5089 255
rect -5097 249 -5095 253
rect -5091 249 -5089 253
rect -5097 247 -5089 249
rect -5097 243 -5095 247
rect -5091 243 -5089 247
rect -5097 241 -5089 243
rect -5097 237 -5095 241
rect -5091 237 -5089 241
rect -5097 235 -5089 237
rect -5097 231 -5095 235
rect -5091 231 -5089 235
rect -5097 230 -5089 231
rect -5097 226 -5095 230
rect -5091 226 -5089 230
rect -5097 224 -5089 226
rect -5097 220 -5095 224
rect -5091 220 -5089 224
rect -5202 218 -5089 220
rect -5202 214 -5195 218
rect -5191 214 -5138 218
rect -5134 214 -5133 218
rect -5129 214 -5126 218
rect -5122 214 -5119 218
rect -5115 214 -5111 218
rect -5107 214 -5105 218
rect -5101 214 -5100 218
rect -5096 214 -5089 218
rect -5202 212 -5089 214
rect -5202 211 -5194 212
rect -5202 207 -5200 211
rect -5196 207 -5194 211
rect -5202 205 -5194 207
rect -5202 201 -5200 205
rect -5196 201 -5194 205
rect -5202 199 -5194 201
rect -5202 195 -5200 199
rect -5196 195 -5194 199
rect -5202 193 -5194 195
rect -5202 189 -5200 193
rect -5196 189 -5194 193
rect -5202 187 -5194 189
rect -5202 183 -5200 187
rect -5196 183 -5194 187
rect -5202 179 -5194 183
rect -5202 175 -5200 179
rect -5196 175 -5194 179
rect -5202 172 -5194 175
rect -5202 168 -5200 172
rect -5196 168 -5194 172
rect -5202 165 -5194 168
rect -5202 161 -5200 165
rect -5196 161 -5194 165
rect -5202 157 -5194 161
rect -5202 153 -5200 157
rect -5196 153 -5194 157
rect -5202 147 -5194 153
rect -5202 143 -5200 147
rect -5196 143 -5194 147
rect -5202 138 -5194 143
rect -5202 134 -5200 138
rect -5196 134 -5194 138
rect -5202 129 -5194 134
rect -5202 125 -5200 129
rect -5196 125 -5194 129
rect -5282 123 -5194 125
rect -5282 119 -5273 123
rect -5269 119 -5266 123
rect -5262 119 -5259 123
rect -5255 119 -5251 123
rect -5247 119 -5245 123
rect -5241 119 -5237 123
rect -5233 119 -5231 123
rect -5227 119 -5223 123
rect -5219 119 -5216 123
rect -5212 119 -5209 123
rect -5205 119 -5204 123
rect -5200 119 -5194 123
rect -5282 118 -5194 119
rect -5282 114 -5280 118
rect -5276 117 -5194 118
rect -5276 114 -5274 117
rect -5282 111 -5274 114
rect -5282 107 -5280 111
rect -5276 107 -5274 111
rect -5282 105 -5274 107
rect -5282 101 -5280 105
rect -5276 101 -5274 105
rect -5282 97 -5274 101
rect -4868 290 -4860 292
rect -4868 286 -4866 290
rect -4862 286 -4860 290
rect -4868 284 -4860 286
rect -4868 280 -4866 284
rect -4862 280 -4860 284
rect -4868 278 -4860 280
rect -4868 274 -4866 278
rect -4862 274 -4860 278
rect -4868 272 -4860 274
rect -4868 268 -4866 272
rect -4862 268 -4860 272
rect -4868 266 -4860 268
rect -4868 262 -4866 266
rect -4862 262 -4860 266
rect -4868 260 -4860 262
rect -4868 256 -4866 260
rect -4862 256 -4860 260
rect -4868 254 -4860 256
rect -4868 250 -4866 254
rect -4862 250 -4860 254
rect -4868 248 -4860 250
rect -4868 244 -4866 248
rect -4862 244 -4860 248
rect -4868 242 -4860 244
rect -4868 238 -4866 242
rect -4862 238 -4860 242
rect -4868 236 -4860 238
rect -4868 232 -4866 236
rect -4862 232 -4860 236
rect -4868 230 -4860 232
rect -4868 226 -4866 230
rect -4862 226 -4860 230
rect -4868 224 -4860 226
rect -4868 220 -4866 224
rect -4862 220 -4860 224
rect -4868 218 -4860 220
rect -4868 214 -4866 218
rect -4862 214 -4860 218
rect -4868 212 -4860 214
rect -4868 208 -4866 212
rect -4862 208 -4860 212
rect -4868 206 -4860 208
rect -4868 202 -4866 206
rect -4862 202 -4860 206
rect -4868 200 -4860 202
rect -4868 196 -4866 200
rect -4862 196 -4860 200
rect -4868 194 -4860 196
rect -4868 190 -4866 194
rect -4862 190 -4860 194
rect -4868 188 -4860 190
rect -4868 184 -4866 188
rect -4862 184 -4860 188
rect -4868 182 -4860 184
rect -4868 178 -4866 182
rect -4862 178 -4860 182
rect -4868 176 -4860 178
rect -4868 172 -4866 176
rect -4862 172 -4860 176
rect -4868 170 -4860 172
rect -4868 166 -4866 170
rect -4862 166 -4860 170
rect -4868 164 -4860 166
rect -4868 160 -4866 164
rect -4862 160 -4860 164
rect -4868 158 -4860 160
rect -4868 154 -4866 158
rect -4862 154 -4860 158
rect -4868 152 -4860 154
rect -4868 148 -4866 152
rect -4862 148 -4860 152
rect -4868 146 -4860 148
rect -4868 142 -4866 146
rect -4862 142 -4860 146
rect -4868 140 -4860 142
rect -4868 136 -4866 140
rect -4862 136 -4860 140
rect -4868 134 -4860 136
rect -4868 130 -4866 134
rect -4862 130 -4860 134
rect -4868 128 -4860 130
rect -4868 124 -4866 128
rect -4862 124 -4860 128
rect -4868 122 -4860 124
rect -4868 118 -4866 122
rect -4862 118 -4860 122
rect -4868 116 -4860 118
rect -4868 112 -4866 116
rect -4862 112 -4860 116
rect -4868 110 -4860 112
rect -4868 106 -4866 110
rect -4862 106 -4860 110
rect -4868 104 -4860 106
rect -4868 100 -4866 104
rect -4862 100 -4860 104
rect -4868 98 -4860 100
rect -4868 94 -4866 98
rect -4862 94 -4860 98
rect -4868 92 -4860 94
rect -4868 88 -4866 92
rect -4862 88 -4860 92
rect -4868 84 -4860 88
<< psubstratepcontact >>
rect -5105 328 -5101 332
rect -5099 328 -5095 332
rect -5093 328 -5089 332
rect -5087 328 -5083 332
rect -5081 328 -5077 332
rect -5073 328 -5069 332
rect -5067 328 -5063 332
rect -5061 328 -5057 332
rect -5055 328 -5051 332
rect -5049 328 -5045 332
rect -5043 328 -5039 332
rect -5037 328 -5033 332
rect -5031 328 -5027 332
rect -5025 328 -5021 332
rect -5019 328 -5015 332
rect -5013 328 -5009 332
rect -5007 328 -5003 332
rect -4999 328 -4995 332
rect -4993 328 -4989 332
rect -4987 328 -4983 332
rect -4981 328 -4977 332
rect -4975 328 -4971 332
rect -4969 328 -4965 332
rect -4963 328 -4959 332
rect -4957 328 -4953 332
rect -4951 328 -4947 332
rect -4945 328 -4941 332
rect -4939 328 -4935 332
rect -4933 328 -4929 332
rect -4925 328 -4921 332
rect -4919 328 -4915 332
rect -4913 328 -4909 332
rect -4907 328 -4903 332
rect -4901 328 -4897 332
rect -4895 328 -4891 332
rect -4889 328 -4885 332
rect -4883 328 -4879 332
rect -4877 328 -4873 332
rect -4871 328 -4867 332
rect -4865 328 -4861 332
rect -4859 328 -4855 332
rect -5114 323 -5110 327
rect -4851 322 -4847 326
rect -5114 316 -5110 320
rect -5114 308 -5110 312
rect -5114 301 -5110 305
rect -5114 295 -5110 299
rect -5114 288 -5110 292
rect -5114 283 -5110 287
rect -5114 278 -5110 282
rect -5114 273 -5110 277
rect -5114 267 -5110 271
rect -5114 261 -5110 265
rect -5114 256 -5110 260
rect -5114 250 -5110 254
rect -5114 244 -5110 248
rect -5114 239 -5110 243
rect -5211 233 -5207 237
rect -5205 233 -5201 237
rect -5199 233 -5195 237
rect -5194 233 -5190 237
rect -5139 233 -5135 237
rect -5134 233 -5130 237
rect -5129 233 -5125 237
rect -5122 233 -5118 237
rect -5217 226 -5213 230
rect -5217 219 -5213 223
rect -5217 214 -5213 218
rect -5217 206 -5213 210
rect -5217 201 -5213 205
rect -5217 196 -5213 200
rect -5217 188 -5213 192
rect -5217 180 -5213 184
rect -5217 173 -5213 177
rect -5217 167 -5213 171
rect -5217 162 -5213 166
rect -5217 154 -5213 158
rect -5217 149 -5213 153
rect -5217 141 -5213 145
rect -5289 136 -5285 140
rect -5283 136 -5279 140
rect -5276 136 -5272 140
rect -5269 136 -5265 140
rect -5262 136 -5258 140
rect -5255 136 -5251 140
rect -5250 136 -5246 140
rect -5245 136 -5241 140
rect -5239 136 -5235 140
rect -5233 136 -5229 140
rect -5227 136 -5223 140
rect -5222 136 -5218 140
rect -5295 128 -5291 132
rect -5295 120 -5291 124
rect -5295 112 -5291 116
rect -5295 105 -5291 109
rect -5295 100 -5291 104
rect -5295 95 -5291 99
rect -5295 89 -5291 93
rect -5295 82 -5291 86
rect -4851 317 -4847 321
rect -4851 311 -4847 315
rect -4851 305 -4847 309
rect -4851 299 -4847 303
rect -4851 293 -4847 297
rect -4851 287 -4847 291
rect -4851 281 -4847 285
rect -4851 275 -4847 279
rect -4851 269 -4847 273
rect -4851 263 -4847 267
rect -4851 257 -4847 261
rect -4851 251 -4847 255
rect -4851 243 -4847 247
rect -4851 237 -4847 241
rect -4851 231 -4847 235
rect -4851 225 -4847 229
rect -4851 219 -4847 223
rect -4851 213 -4847 217
rect -4851 207 -4847 211
rect -4851 201 -4847 205
rect -4851 195 -4847 199
rect -4851 189 -4847 193
rect -4851 183 -4847 187
rect -4851 177 -4847 181
rect -4851 169 -4847 173
rect -4851 163 -4847 167
rect -4851 157 -4847 161
rect -4851 151 -4847 155
rect -4851 145 -4847 149
rect -4851 139 -4847 143
rect -4851 133 -4847 137
rect -4851 127 -4847 131
rect -4851 121 -4847 125
rect -4851 115 -4847 119
rect -4851 109 -4847 113
rect -4851 103 -4847 107
rect -4851 95 -4847 99
rect -4851 89 -4847 93
rect -5295 46 -5291 50
rect -5295 41 -5291 45
rect -4851 83 -4847 87
rect -4851 59 -4847 63
rect -4851 53 -4847 57
rect -5295 33 -5291 37
rect -5295 25 -5291 29
rect -5295 17 -5291 21
rect -5288 10 -5284 14
rect -5281 10 -5277 14
rect -5275 10 -5271 14
rect -5205 10 -5201 14
rect -5197 10 -5193 14
rect -5189 10 -5185 14
rect -5181 10 -5177 14
rect -5173 10 -5169 14
rect -5167 10 -5163 14
rect -5157 10 -5153 14
rect -5149 10 -5145 14
rect -5141 10 -5137 14
rect -5133 10 -5129 14
rect -5124 10 -5120 14
rect -5117 10 -5113 14
rect -5111 10 -5107 14
rect -5106 10 -5102 14
rect -5101 10 -5097 14
rect -5096 10 -5092 14
rect -5091 10 -5087 14
rect -5086 10 -5082 14
rect -5078 10 -5074 14
rect -5069 5 -5065 9
rect -5069 -2 -5065 2
rect -5069 -8 -5065 -4
rect -5069 -13 -5065 -9
rect -5069 -20 -5065 -16
rect -5069 -28 -5065 -24
rect -5069 -35 -5065 -31
rect -5069 -41 -5065 -37
rect -5069 -48 -5065 -44
rect -4851 47 -4847 51
rect -4851 41 -4847 45
rect -4851 35 -4847 39
rect -4851 29 -4847 33
rect -4851 21 -4847 25
rect -4851 15 -4847 19
rect -4851 9 -4847 13
rect -4851 3 -4847 7
rect -4851 -3 -4847 1
rect -4851 -9 -4847 -5
rect -4851 -15 -4847 -11
rect -4851 -21 -4847 -17
rect -4851 -27 -4847 -23
rect -4851 -33 -4847 -29
rect -4851 -39 -4847 -35
rect -4851 -45 -4847 -41
rect -4851 -50 -4847 -46
rect -5069 -55 -5065 -51
rect -4851 -56 -4847 -52
rect -5062 -62 -5058 -58
rect -5056 -62 -5052 -58
rect -5050 -62 -5046 -58
rect -5044 -62 -5040 -58
rect -5038 -62 -5034 -58
rect -5032 -62 -5028 -58
rect -5026 -62 -5022 -58
rect -5020 -62 -5016 -58
rect -5014 -62 -5010 -58
rect -5006 -62 -5002 -58
rect -5000 -62 -4996 -58
rect -4994 -62 -4990 -58
rect -4988 -62 -4984 -58
rect -4982 -62 -4978 -58
rect -4976 -62 -4972 -58
rect -4970 -62 -4966 -58
rect -4964 -62 -4960 -58
rect -4958 -62 -4954 -58
rect -4952 -62 -4948 -58
rect -4946 -62 -4942 -58
rect -4940 -62 -4936 -58
rect -4932 -62 -4928 -58
rect -4926 -62 -4922 -58
rect -4920 -62 -4916 -58
rect -4914 -62 -4910 -58
rect -4908 -62 -4904 -58
rect -4902 -62 -4898 -58
rect -4896 -62 -4892 -58
rect -4890 -62 -4886 -58
rect -4884 -62 -4880 -58
rect -4878 -62 -4874 -58
rect -4872 -62 -4868 -58
rect -4866 -62 -4862 -58
rect -4861 -62 -4857 -58
rect -4856 -62 -4852 -58
<< nsubstratencontact >>
rect -5088 314 -5084 318
rect -5083 314 -5079 318
rect -5078 314 -5074 318
rect -5072 314 -5068 318
rect -5066 314 -5062 318
rect -5058 314 -5054 318
rect -5052 314 -5048 318
rect -5046 314 -5042 318
rect -5040 314 -5036 318
rect -5034 314 -5030 318
rect -5028 314 -5024 318
rect -5022 314 -5018 318
rect -5016 314 -5012 318
rect -5010 314 -5006 318
rect -5004 314 -5000 318
rect -4998 314 -4994 318
rect -4992 314 -4988 318
rect -4986 314 -4982 318
rect -4980 314 -4976 318
rect -4974 314 -4970 318
rect -4968 314 -4964 318
rect -4962 314 -4958 318
rect -4956 314 -4952 318
rect -4950 314 -4946 318
rect -4944 314 -4940 318
rect -4938 314 -4934 318
rect -4932 314 -4928 318
rect -4926 314 -4922 318
rect -4920 314 -4916 318
rect -4914 314 -4910 318
rect -4908 314 -4904 318
rect -4902 314 -4898 318
rect -4896 314 -4892 318
rect -4890 314 -4886 318
rect -4884 314 -4880 318
rect -4878 314 -4874 318
rect -4872 314 -4868 318
rect -5095 309 -5091 313
rect -5095 303 -5091 307
rect -5095 297 -5091 301
rect -4866 310 -4862 314
rect -4866 304 -4862 308
rect -4866 298 -4862 302
rect -5095 291 -5091 295
rect -4866 292 -4862 296
rect -5095 285 -5091 289
rect -5095 277 -5091 281
rect -5095 271 -5091 275
rect -5095 263 -5091 267
rect -5095 255 -5091 259
rect -5095 249 -5091 253
rect -5095 243 -5091 247
rect -5095 237 -5091 241
rect -5095 231 -5091 235
rect -5095 226 -5091 230
rect -5095 220 -5091 224
rect -5195 214 -5191 218
rect -5138 214 -5134 218
rect -5133 214 -5129 218
rect -5126 214 -5122 218
rect -5119 214 -5115 218
rect -5111 214 -5107 218
rect -5105 214 -5101 218
rect -5100 214 -5096 218
rect -5200 207 -5196 211
rect -5200 201 -5196 205
rect -5200 195 -5196 199
rect -5200 189 -5196 193
rect -5200 183 -5196 187
rect -5200 175 -5196 179
rect -5200 168 -5196 172
rect -5200 161 -5196 165
rect -5200 153 -5196 157
rect -5200 143 -5196 147
rect -5200 134 -5196 138
rect -5200 125 -5196 129
rect -5273 119 -5269 123
rect -5266 119 -5262 123
rect -5259 119 -5255 123
rect -5251 119 -5247 123
rect -5245 119 -5241 123
rect -5237 119 -5233 123
rect -5231 119 -5227 123
rect -5223 119 -5219 123
rect -5216 119 -5212 123
rect -5209 119 -5205 123
rect -5204 119 -5200 123
rect -5280 114 -5276 118
rect -5280 107 -5276 111
rect -5280 101 -5276 105
rect -4866 286 -4862 290
rect -4866 280 -4862 284
rect -4866 274 -4862 278
rect -4866 268 -4862 272
rect -4866 262 -4862 266
rect -4866 256 -4862 260
rect -4866 250 -4862 254
rect -4866 244 -4862 248
rect -4866 238 -4862 242
rect -4866 232 -4862 236
rect -4866 226 -4862 230
rect -4866 220 -4862 224
rect -4866 214 -4862 218
rect -4866 208 -4862 212
rect -4866 202 -4862 206
rect -4866 196 -4862 200
rect -4866 190 -4862 194
rect -4866 184 -4862 188
rect -4866 178 -4862 182
rect -4866 172 -4862 176
rect -4866 166 -4862 170
rect -4866 160 -4862 164
rect -4866 154 -4862 158
rect -4866 148 -4862 152
rect -4866 142 -4862 146
rect -4866 136 -4862 140
rect -4866 130 -4862 134
rect -4866 124 -4862 128
rect -4866 118 -4862 122
rect -4866 112 -4862 116
rect -4866 106 -4862 110
rect -4866 100 -4862 104
rect -4866 94 -4862 98
rect -4866 88 -4862 92
<< polysilicon >>
rect -5049 292 -5047 295
rect -5041 292 -5039 295
rect -5033 292 -5031 295
rect -5025 292 -5023 295
rect -5017 292 -5015 295
rect -5009 292 -5007 295
rect -5001 292 -4999 295
rect -4993 292 -4991 295
rect -4985 292 -4983 295
rect -4977 292 -4975 295
rect -4969 292 -4967 295
rect -4961 292 -4959 295
rect -4953 292 -4951 295
rect -4945 292 -4943 295
rect -4937 292 -4935 295
rect -4929 292 -4927 295
rect -4921 292 -4919 295
rect -4913 292 -4911 295
rect -4905 292 -4903 295
rect -4897 292 -4895 295
rect -4889 292 -4887 295
rect -4881 292 -4879 295
rect -5160 146 -5158 149
rect -5136 146 -5134 149
rect -5128 146 -5126 149
rect -5120 146 -5118 149
rect -5112 146 -5110 149
rect -5104 146 -5102 149
rect -5096 146 -5094 149
rect -5088 146 -5086 149
rect -5080 146 -5078 149
rect -5072 146 -5070 149
rect -5258 107 -5256 110
rect -5250 107 -5248 110
rect -5214 101 -5213 103
rect -5258 94 -5256 101
rect -5250 99 -5248 101
rect -5250 97 -5230 99
rect -5258 92 -5249 94
rect -5232 92 -5230 97
rect -5258 86 -5256 89
rect -5239 86 -5237 89
rect -5215 86 -5213 101
rect -5185 98 -5183 101
rect -5258 74 -5256 80
rect -5283 72 -5256 74
rect -5258 66 -5256 72
rect -5239 66 -5237 80
rect -5215 74 -5213 80
rect -5185 74 -5183 92
rect -5160 74 -5158 92
rect -5136 89 -5134 92
rect -5128 89 -5126 92
rect -5120 89 -5118 92
rect -5112 89 -5110 92
rect -5104 89 -5102 92
rect -5096 89 -5094 92
rect -5088 89 -5086 92
rect -5080 89 -5078 92
rect -5072 89 -5070 92
rect -5136 87 -5070 89
rect -5049 89 -5047 92
rect -5041 89 -5039 92
rect -5033 89 -5031 92
rect -5025 89 -5023 92
rect -5017 89 -5015 92
rect -5009 89 -5007 92
rect -5001 89 -4999 92
rect -4993 89 -4991 92
rect -4985 89 -4983 92
rect -4977 89 -4975 92
rect -4969 89 -4967 92
rect -4961 89 -4959 92
rect -4953 89 -4951 92
rect -4945 89 -4943 92
rect -4937 89 -4935 92
rect -4929 89 -4927 92
rect -4921 89 -4919 92
rect -4913 89 -4911 92
rect -4905 89 -4903 92
rect -4897 89 -4895 92
rect -4889 89 -4887 92
rect -4881 89 -4879 92
rect -5049 87 -4878 89
rect -5136 74 -5134 87
rect -5049 74 -5047 87
rect -5214 70 -5213 74
rect -5184 70 -5183 74
rect -5159 70 -5158 74
rect -5135 70 -5134 74
rect -5048 70 -5047 74
rect -5215 66 -5213 70
rect -5258 60 -5256 63
rect -5239 57 -5237 63
rect -5215 60 -5213 63
rect -5283 55 -5237 57
rect -5254 46 -5253 48
rect -5237 46 -5236 48
rect -5185 52 -5183 70
rect -5160 53 -5158 70
rect -5136 58 -5134 70
rect -5049 58 -5047 70
rect -5136 56 -5070 58
rect -5136 53 -5134 56
rect -5128 53 -5126 56
rect -5120 53 -5118 56
rect -5112 53 -5110 56
rect -5104 53 -5102 56
rect -5096 53 -5094 56
rect -5088 53 -5086 56
rect -5080 53 -5078 56
rect -5072 53 -5070 56
rect -5049 56 -4879 58
rect -5049 53 -5047 56
rect -5041 53 -5039 56
rect -5033 53 -5031 56
rect -5025 53 -5023 56
rect -5017 53 -5015 56
rect -5009 53 -5007 56
rect -5001 53 -4999 56
rect -4993 53 -4991 56
rect -4985 53 -4983 56
rect -4977 53 -4975 56
rect -4969 53 -4967 56
rect -4961 53 -4959 56
rect -4953 53 -4951 56
rect -4945 53 -4943 56
rect -4937 53 -4935 56
rect -4929 53 -4927 56
rect -4921 53 -4919 56
rect -4913 53 -4911 56
rect -4905 53 -4903 56
rect -4897 53 -4895 56
rect -4889 53 -4887 56
rect -4881 53 -4879 56
rect -5185 46 -5183 49
rect -5254 37 -5252 46
rect -5237 37 -5235 46
rect -5254 31 -5252 34
rect -5237 31 -5235 34
rect -5160 23 -5158 26
rect -5136 23 -5134 26
rect -5128 23 -5126 26
rect -5120 23 -5118 26
rect -5112 23 -5110 26
rect -5104 23 -5102 26
rect -5096 23 -5094 26
rect -5088 23 -5086 26
rect -5080 23 -5078 26
rect -5072 23 -5070 26
rect -5049 -50 -5047 -47
rect -5041 -50 -5039 -47
rect -5033 -50 -5031 -47
rect -5025 -50 -5023 -47
rect -5017 -50 -5015 -47
rect -5009 -50 -5007 -47
rect -5001 -50 -4999 -47
rect -4993 -50 -4991 -47
rect -4985 -50 -4983 -47
rect -4977 -50 -4975 -47
rect -4969 -50 -4967 -47
rect -4961 -50 -4959 -47
rect -4953 -50 -4951 -47
rect -4945 -50 -4943 -47
rect -4937 -50 -4935 -47
rect -4929 -50 -4927 -47
rect -4921 -50 -4919 -47
rect -4913 -50 -4911 -47
rect -4905 -50 -4903 -47
rect -4897 -50 -4895 -47
rect -4889 -50 -4887 -47
rect -4881 -50 -4879 -47
<< polycontact >>
rect -5218 101 -5214 105
rect -5251 88 -5247 92
rect -5232 88 -5228 92
rect -5287 72 -5283 76
rect -5218 70 -5214 74
rect -5188 70 -5184 74
rect -5163 70 -5159 74
rect -5139 70 -5135 74
rect -5052 70 -5048 74
rect -5287 55 -5283 59
rect -5253 46 -5249 50
rect -5236 46 -5232 50
<< metal1 >>
rect -5115 332 -4846 333
rect -5115 328 -5105 332
rect -5101 328 -5099 332
rect -5095 328 -5093 332
rect -5089 328 -5087 332
rect -5083 328 -5081 332
rect -5077 328 -5073 332
rect -5069 328 -5067 332
rect -5063 328 -5061 332
rect -5057 328 -5055 332
rect -5051 328 -5049 332
rect -5045 328 -5043 332
rect -5039 328 -5037 332
rect -5033 328 -5031 332
rect -5027 328 -5025 332
rect -5021 328 -5019 332
rect -5015 328 -5013 332
rect -5009 328 -5007 332
rect -5003 328 -4999 332
rect -4995 328 -4993 332
rect -4989 328 -4987 332
rect -4983 328 -4981 332
rect -4977 328 -4975 332
rect -4971 328 -4969 332
rect -4965 328 -4963 332
rect -4959 328 -4957 332
rect -4953 328 -4951 332
rect -4947 328 -4945 332
rect -4941 328 -4939 332
rect -4935 328 -4933 332
rect -4929 328 -4925 332
rect -4921 328 -4919 332
rect -4915 328 -4913 332
rect -4909 328 -4907 332
rect -4903 328 -4901 332
rect -4897 328 -4895 332
rect -4891 328 -4889 332
rect -4885 328 -4883 332
rect -4879 328 -4877 332
rect -4873 328 -4871 332
rect -4867 328 -4865 332
rect -4861 328 -4859 332
rect -4855 328 -4846 332
rect -5115 327 -4846 328
rect -5115 323 -5114 327
rect -5110 323 -5109 327
rect -5115 320 -5109 323
rect -5115 316 -5114 320
rect -5110 316 -5109 320
rect -4852 326 -4846 327
rect -4852 322 -4851 326
rect -4847 322 -4846 326
rect -4852 321 -4846 322
rect -5115 312 -5109 316
rect -5115 308 -5114 312
rect -5110 308 -5109 312
rect -5115 305 -5109 308
rect -5115 301 -5114 305
rect -5110 301 -5109 305
rect -5115 299 -5109 301
rect -5115 295 -5114 299
rect -5110 295 -5109 299
rect -5115 292 -5109 295
rect -5115 288 -5114 292
rect -5110 288 -5109 292
rect -5115 287 -5109 288
rect -5115 283 -5114 287
rect -5110 283 -5109 287
rect -5115 282 -5109 283
rect -5115 278 -5114 282
rect -5110 278 -5109 282
rect -5115 277 -5109 278
rect -5115 273 -5114 277
rect -5110 273 -5109 277
rect -5115 271 -5109 273
rect -5115 267 -5114 271
rect -5110 267 -5109 271
rect -5115 265 -5109 267
rect -5115 261 -5114 265
rect -5110 261 -5109 265
rect -5115 260 -5109 261
rect -5115 256 -5114 260
rect -5110 256 -5109 260
rect -5115 254 -5109 256
rect -5115 250 -5114 254
rect -5110 250 -5109 254
rect -5115 248 -5109 250
rect -5190 238 -5140 241
rect -5115 244 -5114 248
rect -5110 244 -5109 248
rect -5115 243 -5109 244
rect -5115 239 -5114 243
rect -5110 239 -5109 243
rect -5115 238 -5109 239
rect -5218 237 -5109 238
rect -5218 233 -5211 237
rect -5207 233 -5205 237
rect -5201 233 -5199 237
rect -5195 233 -5194 237
rect -5190 233 -5139 237
rect -5135 233 -5134 237
rect -5130 233 -5129 237
rect -5125 233 -5122 237
rect -5118 233 -5109 237
rect -5218 232 -5109 233
rect -5096 318 -4861 319
rect -5096 314 -5088 318
rect -5084 314 -5083 318
rect -5079 314 -5078 318
rect -5074 314 -5072 318
rect -5068 314 -5066 318
rect -5062 314 -5058 318
rect -5054 314 -5052 318
rect -5048 314 -5046 318
rect -5042 314 -5040 318
rect -5036 314 -5034 318
rect -5030 314 -5028 318
rect -5024 314 -5022 318
rect -5018 314 -5016 318
rect -5012 314 -5010 318
rect -5006 314 -5004 318
rect -5000 314 -4998 318
rect -4994 314 -4992 318
rect -4988 314 -4986 318
rect -4982 314 -4980 318
rect -4976 314 -4974 318
rect -4970 314 -4968 318
rect -4964 314 -4962 318
rect -4958 314 -4956 318
rect -4952 314 -4950 318
rect -4946 314 -4944 318
rect -4940 314 -4938 318
rect -4934 314 -4932 318
rect -4928 314 -4926 318
rect -4922 314 -4920 318
rect -4916 314 -4914 318
rect -4910 314 -4908 318
rect -4904 314 -4902 318
rect -4898 314 -4896 318
rect -4892 314 -4890 318
rect -4886 314 -4884 318
rect -4880 314 -4878 318
rect -4874 314 -4872 318
rect -4868 314 -4861 318
rect -5096 313 -4866 314
rect -5096 309 -5095 313
rect -5091 309 -5090 313
rect -4867 310 -4866 313
rect -4862 310 -4861 314
rect -5096 307 -5090 309
rect -5096 303 -5095 307
rect -5091 303 -5090 307
rect -5096 301 -5090 303
rect -5096 297 -5095 301
rect -5091 297 -5090 301
rect -5096 295 -5090 297
rect -5096 291 -5095 295
rect -5091 291 -5090 295
rect -5096 289 -5090 291
rect -5096 285 -5095 289
rect -5091 285 -5090 289
rect -5096 281 -5090 285
rect -5096 277 -5095 281
rect -5091 277 -5090 281
rect -5096 275 -5090 277
rect -5096 271 -5095 275
rect -5091 271 -5090 275
rect -5096 267 -5090 271
rect -5096 263 -5095 267
rect -5091 263 -5090 267
rect -5096 259 -5090 263
rect -5096 255 -5095 259
rect -5091 255 -5090 259
rect -5096 253 -5090 255
rect -5096 249 -5095 253
rect -5091 249 -5090 253
rect -5096 247 -5090 249
rect -5096 243 -5095 247
rect -5091 243 -5090 247
rect -5096 241 -5090 243
rect -5096 237 -5095 241
rect -5091 237 -5090 241
rect -5096 235 -5090 237
rect -5218 230 -5212 232
rect -5218 226 -5217 230
rect -5213 226 -5212 230
rect -5218 223 -5212 226
rect -5218 219 -5217 223
rect -5213 219 -5212 223
rect -5190 219 -5140 232
rect -5096 231 -5095 235
rect -5091 231 -5090 235
rect -5096 230 -5090 231
rect -5096 226 -5095 230
rect -5091 226 -5090 230
rect -5096 224 -5090 226
rect -5096 220 -5095 224
rect -5091 220 -5090 224
rect -5096 219 -5090 220
rect -5218 218 -5212 219
rect -5218 214 -5217 218
rect -5213 214 -5212 218
rect -5218 210 -5212 214
rect -5218 206 -5217 210
rect -5213 206 -5212 210
rect -5218 205 -5212 206
rect -5218 201 -5217 205
rect -5213 201 -5212 205
rect -5218 200 -5212 201
rect -5218 196 -5217 200
rect -5213 196 -5212 200
rect -5218 192 -5212 196
rect -5218 188 -5217 192
rect -5213 188 -5212 192
rect -5218 184 -5212 188
rect -5218 180 -5217 184
rect -5213 180 -5212 184
rect -5218 177 -5212 180
rect -5218 173 -5217 177
rect -5213 173 -5212 177
rect -5218 171 -5212 173
rect -5218 167 -5217 171
rect -5213 167 -5212 171
rect -5218 166 -5212 167
rect -5218 162 -5217 166
rect -5213 162 -5212 166
rect -5218 158 -5212 162
rect -5218 154 -5217 158
rect -5213 154 -5212 158
rect -5218 153 -5212 154
rect -5218 149 -5217 153
rect -5213 149 -5212 153
rect -5218 145 -5212 149
rect -5218 141 -5217 145
rect -5213 141 -5212 145
rect -5296 140 -5212 141
rect -5296 136 -5289 140
rect -5285 136 -5283 140
rect -5279 136 -5276 140
rect -5272 136 -5269 140
rect -5265 136 -5262 140
rect -5258 136 -5255 140
rect -5251 136 -5250 140
rect -5246 136 -5245 140
rect -5241 136 -5239 140
rect -5235 136 -5233 140
rect -5229 136 -5227 140
rect -5223 136 -5222 140
rect -5218 136 -5212 140
rect -5296 135 -5212 136
rect -5201 218 -5090 219
rect -5201 214 -5195 218
rect -5191 214 -5138 218
rect -5134 214 -5133 218
rect -5129 214 -5126 218
rect -5122 214 -5119 218
rect -5115 214 -5111 218
rect -5107 214 -5105 218
rect -5101 214 -5100 218
rect -5096 214 -5090 218
rect -5201 213 -5090 214
rect -5080 297 -4882 310
rect -5201 211 -5195 213
rect -5201 207 -5200 211
rect -5196 207 -5195 211
rect -5201 205 -5195 207
rect -5201 201 -5200 205
rect -5196 201 -5195 205
rect -5201 199 -5195 201
rect -5201 195 -5200 199
rect -5196 195 -5195 199
rect -5201 193 -5195 195
rect -5201 189 -5200 193
rect -5196 189 -5195 193
rect -5201 187 -5195 189
rect -5201 183 -5200 187
rect -5196 183 -5195 187
rect -5201 179 -5195 183
rect -5201 175 -5200 179
rect -5196 175 -5195 179
rect -5201 172 -5195 175
rect -5201 168 -5200 172
rect -5196 168 -5195 172
rect -5201 165 -5195 168
rect -5201 161 -5200 165
rect -5196 161 -5195 165
rect -5201 157 -5195 161
rect -5201 153 -5200 157
rect -5196 153 -5195 157
rect -5201 147 -5195 153
rect -5201 143 -5200 147
rect -5196 143 -5195 147
rect -5201 138 -5195 143
rect -5296 132 -5290 135
rect -5296 128 -5295 132
rect -5291 128 -5290 132
rect -5296 124 -5290 128
rect -5201 134 -5200 138
rect -5196 134 -5195 138
rect -5201 129 -5195 134
rect -5201 125 -5200 129
rect -5196 125 -5195 129
rect -5201 124 -5195 125
rect -5296 120 -5295 124
rect -5291 120 -5290 124
rect -5296 116 -5290 120
rect -5296 112 -5295 116
rect -5291 112 -5290 116
rect -5296 109 -5290 112
rect -5296 105 -5295 109
rect -5291 105 -5290 109
rect -5296 104 -5290 105
rect -5296 100 -5295 104
rect -5291 100 -5290 104
rect -5296 99 -5290 100
rect -5296 95 -5295 99
rect -5291 95 -5290 99
rect -5281 123 -5195 124
rect -5281 119 -5273 123
rect -5269 119 -5266 123
rect -5262 119 -5259 123
rect -5255 119 -5251 123
rect -5247 119 -5245 123
rect -5241 119 -5237 123
rect -5233 119 -5231 123
rect -5227 119 -5223 123
rect -5219 119 -5216 123
rect -5212 119 -5209 123
rect -5205 119 -5204 123
rect -5200 119 -5195 123
rect -5281 118 -5195 119
rect -5190 203 -5140 213
rect -5080 203 -5065 297
rect -5046 292 -5042 297
rect -5030 292 -5026 297
rect -5014 292 -5010 297
rect -4998 292 -4994 297
rect -4982 292 -4978 297
rect -4966 292 -4962 297
rect -4950 292 -4946 297
rect -4934 292 -4930 297
rect -4918 292 -4914 297
rect -4902 292 -4898 297
rect -4886 292 -4882 297
rect -4867 308 -4861 310
rect -4867 304 -4866 308
rect -4862 304 -4861 308
rect -4867 302 -4861 304
rect -4867 298 -4866 302
rect -4862 298 -4861 302
rect -4867 296 -4861 298
rect -4867 292 -4866 296
rect -4862 292 -4861 296
rect -5190 153 -5065 203
rect -5281 114 -5280 118
rect -5276 114 -5275 118
rect -5190 115 -5186 153
rect -5281 111 -5275 114
rect -5281 107 -5280 111
rect -5276 107 -5275 111
rect -5281 105 -5275 107
rect -5281 101 -5280 105
rect -5276 101 -5275 105
rect -5281 98 -5275 101
rect -5263 111 -5186 115
rect -5263 107 -5259 111
rect -5243 101 -5218 104
rect -5263 98 -5259 101
rect -5190 98 -5186 111
rect -5165 146 -5161 153
rect -5133 152 -5065 153
rect -5133 146 -5129 152
rect -5117 146 -5113 152
rect -5101 146 -5097 152
rect -5085 146 -5081 152
rect -5069 146 -5065 152
rect -5296 93 -5290 95
rect -5296 89 -5295 93
rect -5291 89 -5290 93
rect -5296 86 -5290 89
rect -5296 82 -5295 86
rect -5291 82 -5290 86
rect -5296 79 -5290 82
rect -5263 95 -5216 98
rect -5263 86 -5259 95
rect -5254 86 -5251 91
rect -5243 86 -5240 95
rect -5235 86 -5232 91
rect -5219 86 -5216 95
rect -5297 72 -5287 75
rect -5254 67 -5251 80
rect -5235 67 -5232 80
rect -5211 74 -5208 80
rect -5181 74 -5178 92
rect -5156 74 -5153 92
rect -5141 86 -5137 92
rect -5125 86 -5121 92
rect -5109 86 -5105 92
rect -5093 86 -5089 92
rect -5077 86 -5073 92
rect -5141 83 -5073 86
rect -5054 86 -5050 92
rect -5038 86 -5034 92
rect -5022 86 -5018 92
rect -5006 86 -5002 92
rect -4990 86 -4986 92
rect -4974 86 -4970 92
rect -4958 86 -4954 92
rect -4942 86 -4938 92
rect -4926 86 -4922 92
rect -4910 86 -4906 92
rect -4894 86 -4890 92
rect -4878 86 -4874 92
rect -5054 83 -4874 86
rect -4867 290 -4861 292
rect -4867 286 -4866 290
rect -4862 286 -4861 290
rect -4867 284 -4861 286
rect -4867 280 -4866 284
rect -4862 280 -4861 284
rect -4867 278 -4861 280
rect -4867 274 -4866 278
rect -4862 274 -4861 278
rect -4867 272 -4861 274
rect -4867 268 -4866 272
rect -4862 268 -4861 272
rect -4867 266 -4861 268
rect -4867 262 -4866 266
rect -4862 262 -4861 266
rect -4867 260 -4861 262
rect -4867 256 -4866 260
rect -4862 256 -4861 260
rect -4867 254 -4861 256
rect -4867 250 -4866 254
rect -4862 250 -4861 254
rect -4867 248 -4861 250
rect -4867 244 -4866 248
rect -4862 244 -4861 248
rect -4867 242 -4861 244
rect -4867 238 -4866 242
rect -4862 238 -4861 242
rect -4867 236 -4861 238
rect -4867 232 -4866 236
rect -4862 232 -4861 236
rect -4867 230 -4861 232
rect -4867 226 -4866 230
rect -4862 226 -4861 230
rect -4867 224 -4861 226
rect -4867 220 -4866 224
rect -4862 220 -4861 224
rect -4867 218 -4861 220
rect -4867 214 -4866 218
rect -4862 214 -4861 218
rect -4867 212 -4861 214
rect -4867 208 -4866 212
rect -4862 208 -4861 212
rect -4867 206 -4861 208
rect -4867 202 -4866 206
rect -4862 202 -4861 206
rect -4867 200 -4861 202
rect -4867 196 -4866 200
rect -4862 196 -4861 200
rect -4867 194 -4861 196
rect -4867 190 -4866 194
rect -4862 190 -4861 194
rect -4867 188 -4861 190
rect -4867 184 -4866 188
rect -4862 184 -4861 188
rect -4867 182 -4861 184
rect -4867 178 -4866 182
rect -4862 178 -4861 182
rect -4867 176 -4861 178
rect -4867 172 -4866 176
rect -4862 172 -4861 176
rect -4867 170 -4861 172
rect -4867 166 -4866 170
rect -4862 166 -4861 170
rect -4867 164 -4861 166
rect -4867 160 -4866 164
rect -4862 160 -4861 164
rect -4867 158 -4861 160
rect -4867 154 -4866 158
rect -4862 154 -4861 158
rect -4867 152 -4861 154
rect -4867 148 -4866 152
rect -4862 148 -4861 152
rect -4867 146 -4861 148
rect -4867 142 -4866 146
rect -4862 142 -4861 146
rect -4867 140 -4861 142
rect -4867 136 -4866 140
rect -4862 136 -4861 140
rect -4867 134 -4861 136
rect -4867 130 -4866 134
rect -4862 130 -4861 134
rect -4867 128 -4861 130
rect -4867 124 -4866 128
rect -4862 124 -4861 128
rect -4867 122 -4861 124
rect -4867 118 -4866 122
rect -4862 118 -4861 122
rect -4867 116 -4861 118
rect -4867 112 -4866 116
rect -4862 112 -4861 116
rect -4867 110 -4861 112
rect -4867 106 -4866 110
rect -4862 106 -4861 110
rect -4867 104 -4861 106
rect -4867 100 -4866 104
rect -4862 100 -4861 104
rect -4867 98 -4861 100
rect -4867 94 -4866 98
rect -4862 94 -4861 98
rect -4867 92 -4861 94
rect -4867 88 -4866 92
rect -4862 88 -4861 92
rect -4867 85 -4861 88
rect -4852 317 -4851 321
rect -4847 317 -4846 321
rect -4852 315 -4846 317
rect -4852 311 -4851 315
rect -4847 311 -4846 315
rect -4852 309 -4846 311
rect -4852 305 -4851 309
rect -4847 305 -4846 309
rect -4852 303 -4846 305
rect -4852 299 -4851 303
rect -4847 299 -4846 303
rect -4852 297 -4846 299
rect -4852 293 -4851 297
rect -4847 293 -4846 297
rect -4852 291 -4846 293
rect -4852 287 -4851 291
rect -4847 287 -4846 291
rect -4852 285 -4846 287
rect -4852 281 -4851 285
rect -4847 281 -4846 285
rect -4852 279 -4846 281
rect -4852 275 -4851 279
rect -4847 275 -4846 279
rect -4852 273 -4846 275
rect -4852 269 -4851 273
rect -4847 269 -4846 273
rect -4852 267 -4846 269
rect -4852 263 -4851 267
rect -4847 263 -4846 267
rect -4852 261 -4846 263
rect -4852 257 -4851 261
rect -4847 257 -4846 261
rect -4852 255 -4846 257
rect -4852 251 -4851 255
rect -4847 251 -4846 255
rect -4852 247 -4846 251
rect -4852 243 -4851 247
rect -4847 243 -4846 247
rect -4852 241 -4846 243
rect -4852 237 -4851 241
rect -4847 237 -4846 241
rect -4852 235 -4846 237
rect -4852 231 -4851 235
rect -4847 231 -4846 235
rect -4852 229 -4846 231
rect -4852 225 -4851 229
rect -4847 225 -4846 229
rect -4852 223 -4846 225
rect -4852 219 -4851 223
rect -4847 219 -4846 223
rect -4852 217 -4846 219
rect -4852 213 -4851 217
rect -4847 213 -4846 217
rect -4852 211 -4846 213
rect -4852 207 -4851 211
rect -4847 207 -4846 211
rect -4852 205 -4846 207
rect -4852 201 -4851 205
rect -4847 201 -4846 205
rect -4852 199 -4846 201
rect -4852 195 -4851 199
rect -4847 195 -4846 199
rect -4852 193 -4846 195
rect -4852 189 -4851 193
rect -4847 189 -4846 193
rect -4852 187 -4846 189
rect -4852 183 -4851 187
rect -4847 183 -4846 187
rect -4852 181 -4846 183
rect -4852 177 -4851 181
rect -4847 177 -4846 181
rect -4852 173 -4846 177
rect -4852 169 -4851 173
rect -4847 169 -4846 173
rect -4852 167 -4846 169
rect -4852 163 -4851 167
rect -4847 163 -4846 167
rect -4852 161 -4846 163
rect -4852 157 -4851 161
rect -4847 157 -4846 161
rect -4852 155 -4846 157
rect -4852 151 -4851 155
rect -4847 151 -4846 155
rect -4852 149 -4846 151
rect -4852 145 -4851 149
rect -4847 145 -4846 149
rect -4852 143 -4846 145
rect -4852 139 -4851 143
rect -4847 139 -4846 143
rect -4852 137 -4846 139
rect -4852 133 -4851 137
rect -4847 133 -4846 137
rect -4852 131 -4846 133
rect -4852 127 -4851 131
rect -4847 127 -4846 131
rect -4852 125 -4846 127
rect -4852 121 -4851 125
rect -4847 121 -4846 125
rect -4852 119 -4846 121
rect -4852 115 -4851 119
rect -4847 115 -4846 119
rect -4852 113 -4846 115
rect -4852 109 -4851 113
rect -4847 109 -4846 113
rect -4852 107 -4846 109
rect -4852 103 -4851 107
rect -4847 103 -4846 107
rect -4852 99 -4846 103
rect -4852 95 -4851 99
rect -4847 95 -4846 99
rect -4852 93 -4846 95
rect -4852 89 -4851 93
rect -4847 89 -4846 93
rect -4852 87 -4846 89
rect -5077 74 -5073 83
rect -4878 74 -4874 83
rect -4852 83 -4851 87
rect -4847 83 -4846 87
rect -4852 80 -4846 83
rect -5251 63 -5249 67
rect -5297 55 -5287 58
rect -5296 50 -5290 51
rect -5296 46 -5295 50
rect -5291 46 -5290 50
rect -5296 45 -5290 46
rect -5296 41 -5295 45
rect -5291 41 -5290 45
rect -5296 37 -5290 41
rect -5262 37 -5259 63
rect -5252 50 -5249 63
rect -5243 57 -5240 63
rect -5235 50 -5232 63
rect -5226 70 -5218 73
rect -5211 70 -5188 74
rect -5181 70 -5163 74
rect -5156 70 -5139 74
rect -5077 70 -5052 74
rect -4878 70 -4845 74
rect -5226 43 -5223 70
rect -5211 67 -5208 70
rect -5246 40 -5223 43
rect -5246 37 -5243 40
rect -5296 33 -5295 37
rect -5291 33 -5290 37
rect -5296 29 -5290 33
rect -5296 25 -5295 29
rect -5291 25 -5290 29
rect -5296 21 -5290 25
rect -5296 17 -5295 21
rect -5291 17 -5290 21
rect -5296 15 -5290 17
rect -5262 30 -5259 33
rect -5225 30 -5222 33
rect -5219 30 -5216 63
rect -5181 53 -5178 70
rect -5156 53 -5153 70
rect -5077 62 -5073 70
rect -4878 62 -4874 70
rect -5262 21 -5212 30
rect -5189 21 -5186 49
rect -5141 59 -5073 62
rect -5141 53 -5137 59
rect -5125 53 -5121 59
rect -5109 53 -5105 59
rect -5093 53 -5089 59
rect -5077 53 -5073 59
rect -5054 59 -4874 62
rect -5054 53 -5050 59
rect -5038 53 -5034 59
rect -5022 53 -5018 59
rect -5006 53 -5002 59
rect -4990 53 -4986 59
rect -4974 53 -4970 59
rect -4958 53 -4954 59
rect -4942 53 -4938 59
rect -4926 53 -4922 59
rect -4910 53 -4906 59
rect -4894 53 -4890 59
rect -4878 53 -4874 59
rect -5165 21 -5161 26
rect -5133 21 -5129 26
rect -5117 21 -5113 26
rect -5101 21 -5097 26
rect -5085 21 -5081 26
rect -5069 21 -5065 26
rect -5262 18 -5058 21
rect -5296 14 -5267 15
rect -5296 10 -5288 14
rect -5284 10 -5281 14
rect -5277 10 -5275 14
rect -5271 10 -5267 14
rect -5296 9 -5267 10
rect -5262 6 -5212 18
rect -5207 14 -5064 15
rect -5207 10 -5205 14
rect -5201 10 -5197 14
rect -5193 10 -5189 14
rect -5185 10 -5181 14
rect -5177 10 -5173 14
rect -5169 10 -5167 14
rect -5163 10 -5157 14
rect -5153 10 -5149 14
rect -5145 10 -5141 14
rect -5137 10 -5133 14
rect -5129 10 -5124 14
rect -5120 10 -5117 14
rect -5113 10 -5111 14
rect -5107 10 -5106 14
rect -5102 10 -5101 14
rect -5097 10 -5096 14
rect -5092 10 -5091 14
rect -5087 10 -5086 14
rect -5082 10 -5078 14
rect -5074 10 -5064 14
rect -5207 9 -5064 10
rect -5070 5 -5069 9
rect -5065 5 -5064 9
rect -5070 2 -5064 5
rect -5070 -2 -5069 2
rect -5065 -2 -5064 2
rect -5070 -4 -5064 -2
rect -5070 -8 -5069 -4
rect -5065 -8 -5064 -4
rect -5070 -9 -5064 -8
rect -5070 -13 -5069 -9
rect -5065 -13 -5064 -9
rect -5070 -16 -5064 -13
rect -5070 -20 -5069 -16
rect -5065 -20 -5064 -16
rect -5070 -24 -5064 -20
rect -5070 -28 -5069 -24
rect -5065 -28 -5064 -24
rect -5070 -31 -5064 -28
rect -5070 -35 -5069 -31
rect -5065 -35 -5064 -31
rect -5070 -37 -5064 -35
rect -5070 -41 -5069 -37
rect -5065 -41 -5064 -37
rect -5070 -44 -5064 -41
rect -5070 -48 -5069 -44
rect -5065 -48 -5064 -44
rect -5070 -51 -5064 -48
rect -5070 -55 -5069 -51
rect -5065 -55 -5064 -51
rect -5061 -51 -5058 18
rect -4852 63 -4846 64
rect -4852 59 -4851 63
rect -4847 59 -4846 63
rect -4852 57 -4846 59
rect -4852 53 -4851 57
rect -4847 53 -4846 57
rect -4852 51 -4846 53
rect -4852 47 -4851 51
rect -4847 47 -4846 51
rect -4852 45 -4846 47
rect -4852 41 -4851 45
rect -4847 41 -4846 45
rect -4852 39 -4846 41
rect -4852 35 -4851 39
rect -4847 35 -4846 39
rect -4852 33 -4846 35
rect -4852 29 -4851 33
rect -4847 29 -4846 33
rect -4852 25 -4846 29
rect -4852 21 -4851 25
rect -4847 21 -4846 25
rect -4852 19 -4846 21
rect -4852 15 -4851 19
rect -4847 15 -4846 19
rect -4852 13 -4846 15
rect -4852 9 -4851 13
rect -4847 9 -4846 13
rect -4852 7 -4846 9
rect -4852 3 -4851 7
rect -4847 3 -4846 7
rect -4852 1 -4846 3
rect -4852 -3 -4851 1
rect -4847 -3 -4846 1
rect -4852 -5 -4846 -3
rect -4852 -9 -4851 -5
rect -4847 -9 -4846 -5
rect -4852 -11 -4846 -9
rect -4852 -15 -4851 -11
rect -4847 -15 -4846 -11
rect -4852 -17 -4846 -15
rect -4852 -21 -4851 -17
rect -4847 -21 -4846 -17
rect -4852 -23 -4846 -21
rect -4852 -27 -4851 -23
rect -4847 -27 -4846 -23
rect -4852 -29 -4846 -27
rect -4852 -33 -4851 -29
rect -4847 -33 -4846 -29
rect -4852 -35 -4846 -33
rect -4852 -39 -4851 -35
rect -4847 -39 -4846 -35
rect -4852 -41 -4846 -39
rect -4852 -45 -4851 -41
rect -4847 -45 -4846 -41
rect -4852 -46 -4846 -45
rect -5046 -51 -5042 -47
rect -5030 -51 -5026 -47
rect -5014 -51 -5010 -47
rect -4998 -51 -4994 -47
rect -4982 -51 -4978 -47
rect -4966 -51 -4962 -47
rect -4950 -51 -4946 -47
rect -4934 -51 -4930 -47
rect -4918 -51 -4914 -47
rect -4902 -51 -4898 -47
rect -4886 -51 -4882 -47
rect -5061 -54 -4882 -51
rect -4852 -50 -4851 -46
rect -4847 -50 -4846 -46
rect -4852 -52 -4846 -50
rect -5070 -57 -5064 -55
rect -4852 -56 -4851 -52
rect -4847 -56 -4846 -52
rect -4852 -57 -4846 -56
rect -5070 -58 -4846 -57
rect -5070 -62 -5062 -58
rect -5058 -62 -5056 -58
rect -5052 -62 -5050 -58
rect -5046 -62 -5044 -58
rect -5040 -62 -5038 -58
rect -5034 -62 -5032 -58
rect -5028 -62 -5026 -58
rect -5022 -62 -5020 -58
rect -5016 -62 -5014 -58
rect -5010 -62 -5006 -58
rect -5002 -62 -5000 -58
rect -4996 -62 -4994 -58
rect -4990 -62 -4988 -58
rect -4984 -62 -4982 -58
rect -4978 -62 -4976 -58
rect -4972 -62 -4970 -58
rect -4966 -62 -4964 -58
rect -4960 -62 -4958 -58
rect -4954 -62 -4952 -58
rect -4948 -62 -4946 -58
rect -4942 -62 -4940 -58
rect -4936 -62 -4932 -58
rect -4928 -62 -4926 -58
rect -4922 -62 -4920 -58
rect -4916 -62 -4914 -58
rect -4910 -62 -4908 -58
rect -4904 -62 -4902 -58
rect -4898 -62 -4896 -58
rect -4892 -62 -4890 -58
rect -4886 -62 -4884 -58
rect -4880 -62 -4878 -58
rect -4874 -62 -4872 -58
rect -4868 -62 -4866 -58
rect -4862 -62 -4861 -58
rect -4857 -62 -4856 -58
rect -4852 -62 -4846 -58
rect -5070 -63 -4846 -62
<< m2contact >>
rect -5190 241 -5140 245
rect -5259 53 -5255 57
rect -5244 53 -5240 57
rect -5262 2 -5212 6
<< metal2 >>
rect -5255 53 -5244 56
<< labels >>
rlabel polycontact -5285 57 -5285 57 1 inB
rlabel polycontact -5285 74 -5285 74 1 inA
rlabel metal1 -5239 18 -5239 18 1 vss
rlabel metal1 -4875 72 -4875 72 1 out
rlabel metal1 -5164 192 -5164 192 1 vdd
<< end >>
