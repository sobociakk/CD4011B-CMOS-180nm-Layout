magic
tech scmos
timestamp 1769750295
<< nwell >>
rect 4628 3552 4994 3696
rect 5492 3552 5858 3696
rect 6372 3553 6738 3697
rect 4627 3537 4994 3552
rect 5491 3537 5858 3552
rect 6371 3538 6738 3553
rect 3025 2715 3184 3081
rect 3169 2714 3184 2715
rect 8166 2971 8181 2972
rect 8166 2605 8325 2971
rect 3025 1522 3184 1888
rect 3169 1521 3184 1522
rect 3025 367 3184 733
rect 3169 366 3184 367
rect 8167 -425 8182 -424
rect 3025 -798 3184 -432
rect 8167 -791 8326 -425
rect 3169 -799 3184 -798
rect 4356 -1472 4723 -1457
rect 5489 -1472 5856 -1457
rect 6580 -1472 6947 -1457
rect 4356 -1616 4722 -1472
rect 5489 -1616 5855 -1472
rect 6580 -1615 6946 -1472
rect 6580 -1616 6665 -1615
rect 6873 -1616 6946 -1615
<< ndiffusion >>
rect 4675 3308 4942 3411
rect 5539 3308 5806 3411
rect 6419 3309 6686 3412
rect 3310 2762 3413 3029
rect 7937 2657 8040 2924
rect 3310 1569 3413 1836
rect 3310 414 3413 681
rect 3310 -751 3413 -484
rect 7938 -739 8041 -472
rect 4408 -1331 4675 -1228
rect 5541 -1331 5808 -1228
rect 6632 -1331 6899 -1228
<< pdiffusion >>
rect 4673 3566 4942 3668
rect 5537 3566 5806 3668
rect 6417 3567 6686 3669
rect 3053 2760 3155 3029
rect 8195 2657 8297 2926
rect 3053 1567 3155 1836
rect 3053 412 3155 681
rect 3053 -753 3155 -484
rect 8196 -739 8298 -470
rect 4408 -1588 4677 -1486
rect 5541 -1588 5810 -1486
rect 6632 -1588 6901 -1486
<< ndcontact >>
rect 4659 3308 4675 3411
rect 4942 3308 4958 3411
rect 5523 3308 5539 3411
rect 5806 3308 5822 3411
rect 6403 3309 6419 3412
rect 6686 3309 6702 3412
rect 3310 3029 3413 3045
rect 3310 2746 3413 2762
rect 7937 2924 8040 2940
rect 7937 2641 8040 2657
rect 3310 1836 3413 1852
rect 3310 1553 3413 1569
rect 3310 681 3413 697
rect 3310 398 3413 414
rect 3310 -484 3413 -468
rect 3310 -767 3413 -751
rect 7938 -472 8041 -456
rect 7938 -755 8041 -739
rect 4392 -1331 4408 -1228
rect 4675 -1331 4691 -1228
rect 5525 -1331 5541 -1228
rect 5808 -1331 5824 -1228
rect 6616 -1331 6632 -1228
rect 6899 -1331 6915 -1228
<< pdcontact >>
rect 4658 3566 4673 3668
rect 4942 3566 4957 3668
rect 5522 3566 5537 3668
rect 5806 3566 5821 3668
rect 6402 3567 6417 3669
rect 6686 3567 6701 3669
rect 3053 3029 3155 3044
rect 3053 2745 3155 2760
rect 8195 2926 8297 2941
rect 8195 2642 8297 2657
rect 3053 1836 3155 1851
rect 3053 1552 3155 1567
rect 3053 681 3155 696
rect 3053 397 3155 412
rect 3053 -484 3155 -469
rect 3053 -768 3155 -753
rect 8196 -470 8298 -455
rect 8196 -754 8298 -739
rect 4393 -1588 4408 -1486
rect 4677 -1588 4692 -1486
rect 5526 -1588 5541 -1486
rect 5810 -1588 5825 -1486
rect 6617 -1588 6632 -1486
rect 6901 -1588 6916 -1486
<< psubstratepdiff >>
rect 4655 3277 4674 3298
rect 4949 3277 4968 3298
rect 5519 3277 5538 3298
rect 5813 3277 5832 3298
rect 6399 3278 6418 3299
rect 6693 3278 6712 3299
rect 3423 3036 3444 3055
rect 3423 2742 3444 2761
rect 7906 2925 7927 2944
rect 7906 2631 7927 2650
rect 3423 1843 3444 1862
rect 3423 1549 3444 1568
rect 3423 688 3444 707
rect 3423 394 3444 413
rect 3423 -477 3444 -458
rect 3423 -771 3444 -752
rect 7907 -471 7928 -452
rect 7907 -765 7928 -746
rect 4382 -1218 4401 -1197
rect 4676 -1218 4695 -1197
rect 5515 -1218 5534 -1197
rect 5809 -1218 5828 -1197
rect 6606 -1218 6625 -1197
rect 6900 -1218 6919 -1197
<< nsubstratendiff >>
rect 4653 3672 4676 3691
rect 4941 3672 4966 3691
rect 5517 3672 5540 3691
rect 5805 3672 5830 3691
rect 6397 3673 6420 3692
rect 6685 3673 6710 3692
rect 3030 3028 3049 3053
rect 3030 2740 3049 2763
rect 8301 2923 8320 2946
rect 8301 2633 8320 2658
rect 3030 1835 3049 1860
rect 3030 1547 3049 1570
rect 3030 680 3049 705
rect 3030 392 3049 415
rect 3030 -485 3049 -460
rect 3030 -773 3049 -750
rect 8302 -473 8321 -450
rect 8302 -763 8321 -738
rect 4384 -1611 4409 -1592
rect 4674 -1611 4697 -1592
rect 5517 -1611 5542 -1592
rect 5807 -1611 5830 -1592
rect 6608 -1611 6633 -1592
rect 6898 -1611 6921 -1592
<< psubstratepcontact >>
rect 4633 3277 4655 3426
rect 4674 3277 4949 3298
rect 4968 3277 4990 3426
rect 5497 3277 5519 3426
rect 5538 3277 5813 3298
rect 5832 3277 5854 3426
rect 6377 3278 6399 3427
rect 6418 3278 6693 3299
rect 6712 3278 6734 3427
rect 3295 3055 3444 3077
rect 3423 2761 3444 3036
rect 3295 2720 3444 2742
rect 7906 2944 8055 2966
rect 7906 2650 7927 2925
rect 7906 2609 8055 2631
rect 3295 1862 3444 1884
rect 3423 1568 3444 1843
rect 3295 1527 3444 1549
rect 3295 707 3444 729
rect 3423 413 3444 688
rect 3295 372 3444 394
rect 3295 -458 3444 -436
rect 3423 -752 3444 -477
rect 3295 -793 3444 -771
rect 7907 -452 8056 -430
rect 7907 -746 7928 -471
rect 7907 -787 8056 -765
rect 4360 -1346 4382 -1197
rect 4401 -1218 4676 -1197
rect 4695 -1346 4717 -1197
rect 5493 -1346 5515 -1197
rect 5534 -1218 5809 -1197
rect 5828 -1346 5850 -1197
rect 6584 -1346 6606 -1197
rect 6625 -1218 6900 -1197
rect 6919 -1346 6941 -1197
<< nsubstratencontact >>
rect 4632 3542 4653 3691
rect 4676 3672 4941 3691
rect 4966 3542 4987 3691
rect 5496 3542 5517 3691
rect 5540 3672 5805 3691
rect 5830 3542 5851 3691
rect 6376 3543 6397 3692
rect 6420 3673 6685 3692
rect 6710 3543 6731 3692
rect 3030 3053 3179 3074
rect 3030 2763 3049 3028
rect 3030 2719 3179 2740
rect 8171 2946 8320 2967
rect 8301 2658 8320 2923
rect 8171 2612 8320 2633
rect 3030 1860 3179 1881
rect 3030 1570 3049 1835
rect 3030 1526 3179 1547
rect 3030 705 3179 726
rect 3030 415 3049 680
rect 3030 371 3179 392
rect 3030 -460 3179 -439
rect 3030 -750 3049 -485
rect 3030 -794 3179 -773
rect 8172 -450 8321 -429
rect 8302 -738 8321 -473
rect 8172 -784 8321 -763
rect 4363 -1611 4384 -1462
rect 4409 -1611 4674 -1592
rect 4697 -1611 4718 -1462
rect 5496 -1611 5517 -1462
rect 5542 -1611 5807 -1592
rect 5830 -1611 5851 -1462
rect 6587 -1611 6608 -1462
rect 6633 -1611 6898 -1592
rect 6921 -1611 6942 -1462
<< metal1 >>
rect 4197 4172 4797 4872
rect 5333 4172 5933 4872
rect 6469 4172 7069 4872
rect 4395 4104 4610 4172
rect 5531 4104 5746 4172
rect 6667 4104 6882 4172
rect 4453 3939 4545 4104
rect 4297 3847 4545 3939
rect 5581 3910 5700 4104
rect 6750 3917 6835 4104
rect 5581 3875 6126 3910
rect 4300 3521 4403 3847
rect 5581 3809 6128 3875
rect 6748 3834 7053 3917
rect 4653 3672 4676 3691
rect 4941 3672 4966 3691
rect 4673 3610 4942 3629
rect 4794 3523 4839 3610
rect 5517 3672 5540 3691
rect 5805 3672 5830 3691
rect 5537 3610 5806 3629
rect 5658 3523 5703 3610
rect 4573 3522 5043 3523
rect 5440 3522 5916 3523
rect 6003 3522 6128 3809
rect 6397 3673 6420 3692
rect 6685 3673 6710 3692
rect 6417 3611 6686 3630
rect 6538 3524 6583 3611
rect 6939 3524 7053 3834
rect 4573 3521 5096 3522
rect 4300 3520 5096 3521
rect 4300 3438 5157 3520
rect 4300 3434 5043 3438
rect 4300 3429 4625 3434
rect 4366 3428 4625 3429
rect 4794 3366 4839 3434
rect 4675 3347 4942 3366
rect 4655 3277 4674 3298
rect 4949 3277 4968 3298
rect 1684 2963 2384 3150
rect 2715 3114 3287 3203
rect 5047 3172 5157 3438
rect 5440 3434 6131 3522
rect 5047 3147 5160 3172
rect 5440 3164 5465 3434
rect 5658 3366 5703 3434
rect 5911 3432 6131 3434
rect 6270 3439 7053 3524
rect 6270 3435 6959 3439
rect 5539 3347 5806 3366
rect 5519 3277 5538 3298
rect 5813 3277 5832 3298
rect 6270 3212 6328 3435
rect 6538 3367 6583 3435
rect 6419 3348 6686 3367
rect 6399 3278 6418 3299
rect 6693 3278 6712 3299
rect 1684 2914 2452 2963
rect 2715 2914 2804 3114
rect 3030 3028 3049 3053
rect 1684 2825 2804 2914
rect 1684 2748 2452 2825
rect 1684 2550 2384 2748
rect 3030 2740 3049 2763
rect 3092 2926 3111 3029
rect 3198 2926 3287 3114
rect 3423 3036 3444 3055
rect 3355 2926 3374 3029
rect 3092 2881 3374 2926
rect 3092 2760 3111 2881
rect 3198 2695 3287 2881
rect 3355 2762 3374 2881
rect 5049 2953 5160 3147
rect 4918 2921 5163 2953
rect 4918 2859 4934 2921
rect 5438 2891 5475 3164
rect 6259 2932 6333 3212
rect 8063 3122 8737 3123
rect 8063 3024 8808 3122
rect 5438 2869 6067 2891
rect 3423 2742 3444 2761
rect 3875 2695 3990 2698
rect 3198 2628 3990 2695
rect 3198 2627 3903 2628
rect 3971 2034 3990 2628
rect 3971 2033 4433 2034
rect 4915 2033 4934 2859
rect 5979 2856 6067 2869
rect 5979 2118 6068 2856
rect 6259 2753 6336 2932
rect 7906 2925 7927 2944
rect 6262 2529 6336 2753
rect 7976 2805 7995 2924
rect 8063 2805 8152 3024
rect 8239 2805 8258 2926
rect 7976 2760 8258 2805
rect 7976 2657 7995 2760
rect 7906 2631 7927 2650
rect 8063 2547 8152 2760
rect 8239 2657 8258 2760
rect 8301 2923 8320 2946
rect 8721 2835 8808 3024
rect 9047 2932 9747 3130
rect 8979 2835 9747 2932
rect 8721 2765 9747 2835
rect 8979 2717 9747 2765
rect 8301 2633 8320 2658
rect 6255 2473 6336 2529
rect 6255 2135 6334 2473
rect 7045 2161 7660 2165
rect 8066 2161 8124 2547
rect 9047 2530 9747 2717
rect 7045 2135 8125 2161
rect 6255 2132 6528 2135
rect 6966 2131 7660 2135
rect 7045 2129 7660 2131
rect 5979 2115 6523 2118
rect 5979 2114 6068 2115
rect 3980 2031 4433 2033
rect 1684 1827 2384 2014
rect 2733 1953 3287 2031
rect 4880 2030 4934 2033
rect 4880 2029 4925 2030
rect 1684 1739 2452 1827
rect 2735 1739 2831 1953
rect 3030 1835 3049 1860
rect 1684 1667 2831 1739
rect 1684 1612 2452 1667
rect 1684 1414 2384 1612
rect 3030 1547 3049 1570
rect 3092 1733 3111 1836
rect 3198 1733 3287 1953
rect 3971 2017 3984 2019
rect 3971 2014 4430 2017
rect 3423 1843 3444 1862
rect 3355 1733 3374 1836
rect 3092 1688 3374 1733
rect 3092 1567 3111 1688
rect 3198 1471 3287 1688
rect 3355 1569 3374 1688
rect 3423 1549 3444 1568
rect 3971 1511 3984 2014
rect 3823 1471 3903 1472
rect 3971 1471 3983 1511
rect 3198 1426 3983 1471
rect 3198 1425 3903 1426
rect 9053 1394 9747 1994
rect 1684 691 2384 878
rect 3198 787 3287 791
rect 3195 781 3903 787
rect 3195 770 3913 781
rect 1684 622 2452 691
rect 3030 680 3049 705
rect 1684 620 2784 622
rect 1684 542 2787 620
rect 1684 476 2452 542
rect 1684 278 2384 476
rect 2706 382 2787 542
rect 3030 392 3049 415
rect 3092 578 3111 681
rect 3198 578 3287 770
rect 3423 688 3444 707
rect 3355 578 3374 681
rect 3092 533 3374 578
rect 3092 412 3111 533
rect 2706 335 2786 382
rect 3198 335 3287 533
rect 3355 414 3374 533
rect 3423 394 3444 413
rect 3891 356 3913 770
rect 2703 285 3289 335
rect 3890 316 3913 356
rect 3890 314 3944 316
rect 3890 312 4477 314
rect 3932 311 4477 312
rect 4922 309 5019 314
rect 3892 297 3911 298
rect 3892 294 4484 297
rect 3892 285 3911 294
rect 1684 -445 2384 -258
rect 3893 -339 3911 285
rect 4764 -39 4814 -33
rect 5007 -39 5019 309
rect 5901 309 6154 312
rect 6833 309 7520 318
rect 5901 306 6320 309
rect 5901 302 6154 306
rect 6769 305 7520 309
rect 5901 275 5924 302
rect 6833 301 7520 305
rect 6150 289 6323 292
rect 4762 -82 5021 -39
rect 3198 -378 3911 -339
rect 3198 -380 3903 -378
rect 1684 -542 2452 -445
rect 3030 -485 3049 -460
rect 1684 -618 2777 -542
rect 1684 -660 2452 -618
rect 1684 -858 2384 -660
rect 2715 -840 2775 -618
rect 3030 -773 3049 -750
rect 3092 -587 3111 -484
rect 3198 -587 3287 -380
rect 3423 -477 3444 -458
rect 3355 -587 3374 -484
rect 3092 -632 3374 -587
rect 3092 -753 3111 -632
rect 3198 -840 3287 -632
rect 3355 -751 3374 -632
rect 4764 -739 4814 -82
rect 4764 -752 4815 -739
rect 3423 -771 3444 -752
rect 2715 -904 3288 -840
rect 4382 -1218 4401 -1197
rect 4676 -1218 4695 -1197
rect 4408 -1286 4675 -1267
rect 4511 -1354 4556 -1286
rect 4768 -1354 4815 -752
rect 5901 -900 5925 275
rect 6150 -271 6175 289
rect 6969 -271 7052 -267
rect 6150 -293 7056 -271
rect 6162 -297 7056 -293
rect 5901 -933 5933 -900
rect 5913 -1089 5933 -933
rect 5515 -1218 5534 -1197
rect 5809 -1218 5828 -1197
rect 5541 -1286 5808 -1267
rect 5644 -1354 5689 -1286
rect 5907 -1354 5938 -1089
rect 6606 -1218 6625 -1197
rect 6900 -1218 6919 -1197
rect 6632 -1286 6899 -1267
rect 6735 -1354 6780 -1286
rect 6969 -1354 7052 -297
rect 7466 -348 7519 301
rect 9050 258 9747 858
rect 7466 -396 8158 -348
rect 7466 -397 7519 -396
rect 7907 -471 7928 -452
rect 7977 -591 7996 -472
rect 8064 -591 8153 -396
rect 8240 -591 8259 -470
rect 7977 -636 8259 -591
rect 7977 -739 7996 -636
rect 7907 -765 7928 -746
rect 8064 -840 8153 -636
rect 8240 -739 8259 -636
rect 8302 -473 8321 -450
rect 9047 -476 9747 -278
rect 8979 -560 9747 -476
rect 8723 -567 9747 -560
rect 8669 -645 9747 -567
rect 8302 -763 8321 -738
rect 8669 -840 8774 -645
rect 8979 -691 9747 -645
rect 8064 -849 8774 -840
rect 8065 -877 8774 -849
rect 8065 -940 8772 -877
rect 9047 -878 9747 -691
rect 4163 -1443 4815 -1354
rect 4163 -1744 4246 -1443
rect 4511 -1530 4556 -1443
rect 4768 -1446 4815 -1443
rect 5382 -1441 5938 -1354
rect 6426 -1440 7052 -1354
rect 5382 -1443 5919 -1441
rect 6426 -1443 6977 -1440
rect 4408 -1549 4677 -1530
rect 4384 -1611 4409 -1592
rect 4674 -1611 4697 -1592
rect 4163 -1747 4573 -1744
rect 4163 -1845 4576 -1747
rect 5382 -1752 5487 -1443
rect 5644 -1530 5689 -1443
rect 5541 -1549 5810 -1530
rect 5517 -1611 5542 -1592
rect 5807 -1611 5830 -1592
rect 5382 -1837 5713 -1752
rect 6426 -1770 6539 -1443
rect 6735 -1530 6780 -1443
rect 6632 -1549 6901 -1530
rect 6608 -1611 6633 -1592
rect 6898 -1611 6921 -1592
rect 6426 -1835 6845 -1770
rect 4486 -1972 4576 -1845
rect 5596 -1972 5712 -1837
rect 6732 -1972 6845 -1835
rect 4416 -2040 4631 -1972
rect 5552 -2040 5767 -1972
rect 6688 -2040 6903 -1972
rect 4229 -2740 4829 -2040
rect 5365 -2740 5965 -2040
rect 6501 -2740 7101 -2040
<< m2contact >>
rect 4763 3691 4870 3710
rect 5619 3691 5726 3710
rect 6507 3692 6614 3711
rect 4769 3258 4876 3277
rect 5612 3257 5719 3277
rect 6523 3258 6630 3278
rect 2990 2826 3030 2951
rect 3444 2854 3486 2980
rect 7844 2779 7906 2904
rect 8320 2746 8376 2870
rect 2990 1638 3030 1763
rect 3444 1641 3487 1765
rect 2990 482 3030 607
rect 3444 492 3487 616
rect 2990 -684 3030 -560
rect 3444 -667 3487 -542
rect 4446 -1197 4654 -1171
rect 5608 -1197 5798 -1171
rect 6652 -1197 6860 -1171
rect 7845 -743 7907 -617
rect 8321 -697 8376 -569
rect 4445 -1635 4654 -1611
rect 5572 -1635 5781 -1611
rect 6665 -1635 6873 -1611
<< metal2 >>
rect 4197 4172 4797 4872
rect 5333 4172 5933 4872
rect 6469 4172 7069 4872
rect 2952 3711 8415 3747
rect 2952 3710 6507 3711
rect 2952 3272 2989 3710
rect 6614 3710 8415 3711
rect 3444 3277 4602 3278
rect 6249 3277 6523 3278
rect 2952 3269 2990 3272
rect 1684 2550 2384 3150
rect 1684 1414 2384 2014
rect 1684 278 2384 878
rect 1684 -858 2384 -258
rect 2953 -1634 2990 3269
rect 3444 3258 4769 3277
rect 4876 3274 5043 3277
rect 5286 3274 5612 3277
rect 4876 3258 5612 3274
rect 3444 3257 5612 3258
rect 5719 3258 6523 3277
rect 6630 3258 7906 3278
rect 5719 3257 7906 3258
rect 3444 3231 7906 3257
rect 3444 3105 3495 3231
rect 4534 3229 4585 3231
rect 5033 3230 5336 3231
rect 3444 2980 3496 3105
rect 3486 2854 3496 2980
rect 3444 2585 3496 2854
rect 3444 2040 3497 2585
rect 4535 2204 4585 3229
rect 7836 3082 7906 3231
rect 6628 3041 7906 3082
rect 6628 2921 6681 3041
rect 6628 2904 6683 2921
rect 6630 2305 6683 2904
rect 7836 2904 7906 3041
rect 7836 2779 7844 2904
rect 7836 2099 7906 2779
rect 8376 2744 8415 3710
rect 9047 2530 9747 3130
rect 6558 2060 6608 2062
rect 3444 1765 3496 2040
rect 4463 1958 4513 1961
rect 3487 1641 3496 1765
rect 3444 1526 3496 1641
rect 3444 877 3494 1526
rect 4464 1318 4512 1958
rect 6556 1323 6608 2060
rect 7835 2048 7906 2099
rect 7835 1707 7904 2048
rect 7835 1706 8369 1707
rect 8416 1706 8522 1707
rect 9053 1706 9747 1994
rect 7835 1655 9747 1706
rect 8378 1654 9747 1655
rect 9053 1394 9747 1654
rect 8372 1323 8418 1324
rect 5405 1318 8427 1323
rect 4464 1248 8427 1318
rect 4464 1243 7507 1248
rect 4464 1238 4512 1243
rect 3444 842 4635 877
rect 3444 616 3494 842
rect 4582 652 4633 842
rect 3487 492 3494 616
rect 3444 377 3494 492
rect 4583 484 4633 652
rect 3444 -542 3495 377
rect 4510 123 4562 241
rect 5426 123 5467 1243
rect 7861 686 7904 690
rect 7835 684 7904 686
rect 6427 648 7904 684
rect 6426 613 7904 648
rect 6426 479 6476 613
rect 6354 123 6404 236
rect 4510 84 6404 123
rect 3487 -667 3495 -542
rect 3444 -794 3495 -667
rect 3442 -1150 3495 -794
rect 7835 -340 7904 613
rect 8372 581 8418 1248
rect 9050 581 9747 858
rect 8372 576 9747 581
rect 8378 529 9747 576
rect 8378 149 8413 529
rect 9050 258 9747 529
rect 7835 -617 7905 -340
rect 7835 -743 7845 -617
rect 7835 -868 7905 -743
rect 7836 -989 7905 -868
rect 6979 -1150 7267 -1148
rect 7835 -1150 7906 -989
rect 3442 -1171 7906 -1150
rect 3442 -1194 4446 -1171
rect 3445 -1197 4446 -1194
rect 4654 -1197 5608 -1171
rect 5798 -1197 6652 -1171
rect 6860 -1193 7906 -1171
rect 6860 -1197 6981 -1193
rect 7166 -1197 7906 -1193
rect 3445 -1198 3492 -1197
rect 2953 -1635 3415 -1634
rect 8376 -1635 8415 149
rect 9047 -878 9747 -278
rect 2953 -1673 8415 -1635
rect 4229 -2740 4829 -2040
rect 5365 -2740 5965 -2040
rect 6501 -2740 7101 -2040
<< metal3 >>
rect 4197 4172 4797 4872
rect 5333 4172 5933 4872
rect 6469 4172 7069 4872
rect 1684 2550 2384 3150
rect 9047 2530 9747 3130
rect 1684 1414 2384 2014
rect 9053 1394 9747 1994
rect 1684 278 2384 878
rect 9050 258 9747 858
rect 1684 -858 2384 -258
rect 9047 -878 9747 -278
rect 4229 -2740 4829 -2040
rect 5365 -2740 5965 -2040
rect 6501 -2740 7101 -2040
<< metal4 >>
rect 4197 4172 4797 4872
rect 5333 4172 5933 4872
rect 6469 4172 7069 4872
rect 1684 2550 2384 3150
rect 9047 2530 9747 3130
rect 1684 1414 2384 2014
rect 9053 1394 9747 1994
rect 1684 278 2384 878
rect 9050 258 9747 858
rect 1684 -858 2384 -258
rect 9047 -878 9747 -278
rect 4229 -2740 4829 -2040
rect 5365 -2740 5965 -2040
rect 6501 -2740 7101 -2040
<< m6contact >>
rect 4197 4172 4797 4872
rect 5333 4172 5933 4872
rect 6469 4172 7069 4872
rect 1684 2550 2384 3150
rect 9047 2530 9747 3130
rect 1684 1414 2384 2014
rect 9053 1394 9747 1994
rect 1684 278 2384 878
rect 9050 258 9747 858
rect 1684 -858 2384 -258
rect 9047 -878 9747 -278
rect 4229 -2740 4829 -2040
rect 5365 -2740 5965 -2040
rect 6501 -2740 7101 -2040
<< glass >>
rect 4227 4202 4767 4842
rect 5363 4202 5903 4842
rect 6499 4202 7039 4842
rect 1714 2580 2354 3120
rect 9077 2560 9717 3100
rect 1714 1444 2354 1984
rect 9077 1424 9717 1964
rect 1714 308 2354 848
rect 9077 288 9717 828
rect 1714 -828 2354 -288
rect 9077 -848 9717 -308
rect 4259 -2710 4799 -2070
rect 5395 -2710 5935 -2070
rect 6531 -2710 7071 -2070
use nand  nand_3
timestamp 1769746565
transform 1 0 11820 0 1 2060
box -5297 -64 -4845 334
use nand  nand_2
timestamp 1769746565
transform 1 0 11616 0 1 234
box -5297 -64 -4845 334
use nand  nand_1
timestamp 1769746565
transform 1 0 9773 0 1 239
box -5297 -64 -4845 334
use nand  nand_0
timestamp 1769746565
transform 1 0 9725 0 1 1959
box -5297 -64 -4845 334
<< labels >>
rlabel m6contact 9130 1686 9130 1686 1 vdd
rlabel m6contact 9139 564 9139 564 1 vss
<< end >>
